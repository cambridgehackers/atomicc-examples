`ifndef __configCounter_GENERATED__VH__
`define __configCounter_GENERATED__VH__

//METASTART; ConfigCounter
//METAEXCLUSIVE; decrement__ENA; maybeDecrement
//METAGUARD; decrement; 1;
//METAGUARD; maybeDecrement; 1;
//METAGUARD; increment; 1;
//METAGUARD; read; 1;
//METAGUARD; positive; 1;
//METABEFORE; RULE$react__ENA; :decrement__ENA; :increment__ENA; :maybeDecrement
//METAGUARD; RULE$react; 1;
//METARULES; RULE$react
`endif
