interface P7WrapIfc;
    logic [54 - 1:0] MIO;
endinterface
