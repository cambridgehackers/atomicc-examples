`ifndef __clock_GENERATED__VH__
`define __clock_GENERATED__VH__

//METASTART; ModFt600
//METAINTERNAL; iobufs0; IOBUF;
//METAINTERNAL; iobufs1; IOBUF;
//METAINTERNAL; iobufs2; IOBUF;
//METAINTERNAL; iobufs3; IOBUF;
//METAINTERNAL; iobufs4; IOBUF;
//METAINTERNAL; iobufs5; IOBUF;
//METAINTERNAL; iobufs6; IOBUF;
//METAINTERNAL; iobufs7; IOBUF;
//METAINTERNAL; iobufs8; IOBUF;
//METAINTERNAL; iobufs9; IOBUF;
//METAINTERNAL; iobufs10; IOBUF;
//METAINTERNAL; iobufs11; IOBUF;
//METAINTERNAL; iobufs12; IOBUF;
//METAINTERNAL; iobufs13; IOBUF;
//METAINTERNAL; iobufs14; IOBUF;
//METAINTERNAL; iobufs15; IOBUF;
//METAGUARD; RULE$handshake; 1;
//METAGUARD; RULE$iobufs_0; 1;
//METAGUARD; RULE$iobufs_10; 1;
//METAGUARD; RULE$iobufs_11; 1;
//METAGUARD; RULE$iobufs_12; 1;
//METAGUARD; RULE$iobufs_13; 1;
//METAGUARD; RULE$iobufs_14; 1;
//METAGUARD; RULE$iobufs_15; 1;
//METAGUARD; RULE$iobufs_1; 1;
//METAGUARD; RULE$iobufs_2; 1;
//METAGUARD; RULE$iobufs_3; 1;
//METAGUARD; RULE$iobufs_4; 1;
//METAGUARD; RULE$iobufs_5; 1;
//METAGUARD; RULE$iobufs_6; 1;
//METAGUARD; RULE$iobufs_7; 1;
//METAGUARD; RULE$iobufs_8; 1;
//METAGUARD; RULE$iobufs_9; 1;
//METARULES; RULE$handshake; RULE$iobufs_0; RULE$iobufs_1; RULE$iobufs_10; RULE$iobufs_11; RULE$iobufs_12; RULE$iobufs_13; RULE$iobufs_14; RULE$iobufs_15; RULE$iobufs_2; RULE$iobufs_3; RULE$iobufs_4; RULE$iobufs_5; RULE$iobufs_6; RULE$iobufs_7; RULE$iobufs_8; RULE$iobufs_9
`endif
