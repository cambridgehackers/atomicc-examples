interface I2C_Pins;
    logic  scl;
    logic  sda;
endinterface
