`ifndef __configCounter_GENERATED__VH__
`define __configCounter_GENERATED__VH__

//METASTART; ConfigCounter
//METAEXCLUSIVE; ifc$decrement__ENA; ifc$maybeDecrement
//METAGUARD; ifc$decrement; 1;
//METAGUARD; ifc$maybeDecrement; 1;
//METAGUARD; ifc$increment; 1;
//METAGUARD; ifc$read; 1;
//METAGUARD; ifc$positive; 1;
//METABEFORE; RULE$react__ENA; :ifc$decrement__ENA; :ifc$increment__ENA; :ifc$maybeDecrement
//METAGUARD; RULE$react; 1;
//METARULES; RULE$react
`endif
