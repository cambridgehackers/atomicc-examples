`include "atomicclib.vh"

//METASTART; GrayCounter
//METAINTERNAL; __traceMemory; Trace(width=4,depth=1024,sensitivity=99,head=77);
//METAGUARD; increment; 1'd1;
//METAGUARD; decrement; 1'd1;
//METAGUARD; readGray; 1'd1;
//METAGUARD; writeGray; 1'd1;
//METAGUARD; readBin; 1'd1;
//METAGUARD; writeBin; 1'd1;
//METAGUARD; RULE$incdec; increment__ENA != decrement__ENA;
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$incdec; RULE$init
