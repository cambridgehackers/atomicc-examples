`include "atomicclib.vh"

//METASTART; BusyCtr
//METAEXCLUSIVE; startSignal__ENA; RULE$decRule__ENA
//METAGUARD; startSignal; counter == 0;
//METAGUARD; busy; 1'd1;
//METAGUARD; RULE$decRule; counter != 0;
//METAGUARD; RULE$verify0; 1'd1;
//METARULES; RULE$decRule; RULE$verify0
