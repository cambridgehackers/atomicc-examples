`include "atomicclib.vh"

//METASTART; ConfigCounter
//METAGUARD; decrement; 1'd1;
//METAGUARD; maybeDecrement; 1'd1;
//METAGUARD; increment; 1'd1;
//METAGUARD; read; 1'd1;
//METAGUARD; positive; 1'd1;
//METAGUARD; RULE$react; 1'd1;
//METARULES; RULE$react
