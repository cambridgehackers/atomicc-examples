`include "atomicclib.vh"

//METASTART; P7Wrap
//METAINTERNAL; pps; PS7;
//METAINTERNAL; pclockTop; ClockTop;
//METAINTERNAL; tsda0; IOBUF;
//METAINTERNAL; tscl0; IOBUF;
//METAINTERNAL; tsda1; IOBUF;
//METAINTERNAL; tscl1; IOBUF;
//METAGUARD; MAXIGP0_I.R; 0 != pps$MAXIGP0RREADY;
//METAGUARD; MAXIGP0_I.B; 0 != pps$MAXIGP0BREADY;
//METAGUARD; RULE$init; 1'd1;
//METAINVOKE; RULE$gp0ar__ENA; :MAXIGP0_O.AR__ENA;
//METAGUARD; RULE$gp0ar; pps$MAXIGP0ARVALID && MAXIGP0_O.AR__RDY;
//METAINVOKE; RULE$gp0aw__ENA; :MAXIGP0_O.AW__ENA;
//METAGUARD; RULE$gp0aw; pps$MAXIGP0AWVALID && MAXIGP0_O.AW__RDY;
//METAINVOKE; RULE$gp0w__ENA; :MAXIGP0_O.W__ENA;
//METAGUARD; RULE$gp0w; pps$MAXIGP0WVALID && MAXIGP0_O.W__RDY;
//METARULES; RULE$init; RULE$gp0ar; RULE$gp0aw; RULE$gp0w
//METASTART; ZynqTop
//METAINTERNAL; ps7_ps7_foo; P7Wrap;
//METAINTERNAL; test; AxiTop;
//METAINTERNAL; ps7_fclk_0_c; BUFG;
//METAINTERNAL; ps7_freset_0_r; BUFG;
//METAINTERNAL; bscan; Bscan(id=3,width=32);
//METAGUARD; RULE$init; 1'd1;
//METAEXCLUSIVE; readUser.enq__ENA; RULE$resetOneShot__ENA
//METAGUARD; readUser.enq; 1'd1;
//METAGUARD; RULE$resetOneShot; 0 != resetFunnel;
//METARULES; RULE$init; RULE$resetOneShot
//METACONNECT; test$MAXIGP0_O.AR__ENA; ps7_ps7_foo$MAXIGP0_O.AR__ENA
//METACONNECT; test$MAXIGP0_O.AR__RDY; ps7_ps7_foo$MAXIGP0_O.AR__RDY
//METACONNECT; test$MAXIGP0_O.AW__ENA; ps7_ps7_foo$MAXIGP0_O.AW__ENA
//METACONNECT; test$MAXIGP0_O.AW__RDY; ps7_ps7_foo$MAXIGP0_O.AW__RDY
//METACONNECT; test$MAXIGP0_O.W__ENA; ps7_ps7_foo$MAXIGP0_O.W__ENA
//METACONNECT; test$MAXIGP0_O.W__RDY; ps7_ps7_foo$MAXIGP0_O.W__RDY
//METACONNECT; test$MAXIGP0_I.R__ENA; ps7_ps7_foo$MAXIGP0_I.R__ENA
//METACONNECT; test$MAXIGP0_I.R__RDY; ps7_ps7_foo$MAXIGP0_I.R__RDY
//METACONNECT; test$MAXIGP0_I.B__ENA; ps7_ps7_foo$MAXIGP0_I.B__ENA
//METACONNECT; test$MAXIGP0_I.B__RDY; ps7_ps7_foo$MAXIGP0_I.B__RDY
//METACONNECT; readUser.enq__ENA; bscan$fromBscan.enq__ENA
//METACONNECT; readUser.enq__RDY; bscan$fromBscan.enq__RDY
