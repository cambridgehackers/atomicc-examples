`ifndef __funnel_GENERATED__VH__
`define __funnel_GENERATED__VH__

//METASTART; FunnelHalfBase
//METAGUARD; input$enq; 1;
`endif
