`ifndef __funnel_GENERATED__VH__
`define __funnel_GENERATED__VH__

`endif
