
`define BSV_RESET_VALUE 1'b0
`define MAX_IN_WIDTH 128
`define MAX_OUT_WIDTH 128
`define MAX_BUS_WIDTH 32
`define IfcNames_EchoIndicationH2S  16'd5
`define IfcNames_EchoRequestS2H     16'd6
