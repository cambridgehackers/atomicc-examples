`include "zynqTop.generated.vh"

`default_nettype none
module Fifo1old_OC_22 (input wire CLK, input wire nRST,
    input wire in$enq__ENA,
    input wire [31:0]in$enq$v,
    output wire in$enq__RDY,
    input wire out$deq__ENA,
    output wire out$deq__RDY,
    output wire [31:0]out$first,
    output wire out$first__RDY);
    reg [31:0]element$data;
    reg full;
    Fifo1Base_OC_18 fifo (.CLK(CLK), .nRST(nRST),
        .in$enq__ENA(0),
        .in$enq$v(0),
        .in$enq__RDY(),
        .out$deq__ENA(0),
        .out$deq__RDY(),
        .out$first(),
        .out$first__RDY());
    assign in$enq__RDY = !full;
    assign out$deq__RDY = full;
    assign out$first = { element$data };
    assign out$first__RDY = full;

    always @( posedge CLK) begin
      if (!nRST) begin
        element$data <= 0;
        full <= 0;
      end // nRST
      else begin
        if (in$enq__ENA & ( !full )) begin // in$enq__ENA
            { element$data } <= in$enq$v;
            full <= 1;
        end; // End of in$enq__ENA
        if (out$deq__ENA & full) begin // out$deq__ENA
            full <= 0;
        end; // End of out$deq__ENA
      end
    end // always @ (posedge CLK)
endmodule 

`default_nettype wire    // set back to default value
