`ifndef __fifo_GENERATED__VH__
`define __fifo_GENERATED__VH__

//METASTART; l_module_OC_Fifo1
//METAEXCLUSIVE; out$deq; in$enq
//METAGUARD; out$deq; full;
//METAGUARD; in$enq; full ^ 1;
//METABEFORE; out$first; :in$enq
//METAGUARD; out$first; full;
`endif
