`ifndef __fifo_GENERATED__VH__
`define __fifo_GENERATED__VH__

//METASTART; l_module_OC_Fifo1
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; full  ^ 1;
//METAGUARD; out$deq; 0 != full ;
//METAGUARD; out$first; 0 != full ;
`endif
