`include "rulec.generated.vh"

module CONNECTNET2 (
    input IN1,
    input IN2,
    output OUT1,
    output OUT2);
    wire CLK;
    wire nRST;
    wire assign__ENA;
    assign assign__ENA = 1;
    assign OUT1 = IN1 ;
    assign OUT2 = IN2 ;
endmodule 

