`define TopAppendPort
`define TopAppendCode
