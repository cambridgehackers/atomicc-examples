`include "atomicclib.vh"

//METASTART; Printf
//METAGUARD; enq; 1'd1;
