`ifndef __connectNet2_GENERATED__VH__
`define __connectNet2_GENERATED__VH__
`include "atomicclib.vh"

`ifndef __CNCONNECTNET2_DEF__
`define __CNCONNECTNET2_DEF__
interface CNCONNECTNET2;
    logic  IN1;
    logic  IN2;
    logic  OUT1;
    logic  OUT2;
    modport server (input  IN1, IN2,
                    output OUT1, OUT2);
    modport client (output IN1, IN2,
                    input  OUT1, OUT2);
endinterface
`endif
`ifndef __PipeIn_OC_0_DEF__
`define __PipeIn_OC_0_DEF__
interface PipeIn_OC_0#(dataWidth = 32, funnelWidth = 99);
    logic enq__ENA;
    logic [dataWidth - 1:0] enq$v;
    logic enq__RDY;
    modport server (input  enq__ENA, enq$v,
                    output enq__RDY);
    modport client (output enq__ENA, enq$v,
                    input  enq__RDY);
endinterface
`endif
`ifndef __PipeIn_OC_1_DEF__
`define __PipeIn_OC_1_DEF__
interface PipeIn_OC_1#(dataWidth = 32, funnelWidth = 99);
    logic enq__ENA;
    logic [dataWidth - 1:0] enq$v;
    logic enq__RDY;
    modport server (input  enq__ENA, enq$v,
                    output enq__RDY);
    modport client (output enq__ENA, enq$v,
                    input  enq__RDY);
endinterface
`endif
`ifndef __PipeIn_DEF__
`define __PipeIn_DEF__
interface PipeIn;
    logic enq__ENA;
    logic [(16 + 128) - 1:0] enq$v;
    logic enq__RDY;
    modport server (input  enq__ENA, enq$v,
                    output enq__RDY);
    modport client (output enq__ENA, enq$v,
                    input  enq__RDY);
endinterface
`endif
//METASTART; CONNECTNET2
//METAGUARD; RULE$assign; 1;
//METARULES; RULE$assign
`endif
