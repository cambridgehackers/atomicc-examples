`include "atomicclib.vh"

//METASTART; IobufVec
//METAINTERNAL; iobufs0; IOBUF;
//METAGUARD; RULE$iobufs; 1'd1;
//METARULES; RULE$iobufs
