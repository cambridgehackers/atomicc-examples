`ifndef __gear1toN_GENERATED__VH__
`define __gear1toN_GENERATED__VH__

//METASTART; Gear1toNBase
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; !( c == 4 );
//METAGUARD; out$deq; c == 4;
//METAGUARD; out$first; c == 4;
`endif
