`ifndef __fifo_GENERATED__VH__
`define __fifo_GENERATED__VH__

//METASTART; l_module_OC_Fifo1
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; full  ^ 1;
//METAGUARD; out$deq; full ;
//METAGUARD; out$first; full ;
`endif
