`include "atomicclib.vh"

//METASTART; BRAM
//METAGUARD; write; 1'd1;
//METAGUARD; read; 1'd1;
//METAGUARD; dataOut; afterRead != 0;
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$init
