`include "zynqTop.generated.vh"

module ZynqTop (
    output CLK,
    output nRST,
    output [3:0]FCLKCLK,
    inout DDRA,
    input [3:0]DDRARB,
    inout DDRBA,
    inout DDRCASB,
    inout DDRCKE,
    inout DDRCKN,
    inout DDRCKP,
    inout DDRCSB,
    inout DDRDM,
    inout DDRDQ,
    inout DDRDQSN,
    inout DDRDQSP,
    inout DDRDRSTB,
    inout DDRODT,
    inout DDRRASB,
    inout DDRVRN,
    inout DDRVRP,
    inout DDRWEB,
    input [19:0]IRQF2P,
    output [28:0]IRQP2F,
    inout MIO,
    input MAXIGP0ACLK,
    output [31:0]MAXIGP0ARADDR,
    output [1:0]MAXIGP0ARBURST,
    output [3:0]MAXIGP0ARCACHE,
    output MAXIGP0ARESETN,
    output [11:0]MAXIGP0ARID,
    output [3:0]MAXIGP0ARLEN,
    output [1:0]MAXIGP0ARLOCK,
    output [2:0]MAXIGP0ARPROT,
    output [3:0]MAXIGP0ARQOS,
    input MAXIGP0ARREADY,
    output [1:0]MAXIGP0ARSIZE,
    output MAXIGP0ARVALID,
    output [31:0]MAXIGP0AWADDR,
    output [1:0]MAXIGP0AWBURST,
    output [3:0]MAXIGP0AWCACHE,
    output [11:0]MAXIGP0AWID,
    output [3:0]MAXIGP0AWLEN,
    output [1:0]MAXIGP0AWLOCK,
    output [2:0]MAXIGP0AWPROT,
    output [3:0]MAXIGP0AWQOS,
    input MAXIGP0AWREADY,
    output [1:0]MAXIGP0AWSIZE,
    output MAXIGP0AWVALID,
    input [11:0]MAXIGP0BID,
    output MAXIGP0BREADY,
    input [1:0]MAXIGP0BRESP,
    input MAXIGP0BVALID,
    input [31:0]MAXIGP0RDATA,
    input [11:0]MAXIGP0RID,
    input MAXIGP0RLAST,
    output MAXIGP0RREADY,
    input [1:0]MAXIGP0RRESP,
    input MAXIGP0RVALID,
    output [31:0]MAXIGP0WDATA,
    output [11:0]MAXIGP0WID,
    output MAXIGP0WLAST,
    input MAXIGP0WREADY,
    output [3:0]MAXIGP0WSTRB,
    output MAXIGP0WVALID,
    inout PSCLK,
    inout PSPORB,
    inout PSSRSTB);
    wire init__ENA;
    wire pps$DMA0ACLK;
    wire pps$DMA0DAREADY;
    wire [1:0]pps$DMA0DATYPE;
    wire pps$DMA0DAVALID;
    wire pps$DMA0DRLAST;
    wire pps$DMA0DRREADY;
    wire [1:0]pps$DMA0DRTYPE;
    wire pps$DMA0DRVALID;
    wire pps$DMA0RSTN;
    wire pps$DMA1ACLK;
    wire pps$DMA1DAREADY;
    wire [1:0]pps$DMA1DATYPE;
    wire pps$DMA1DAVALID;
    wire pps$DMA1DRLAST;
    wire pps$DMA1DRREADY;
    wire [1:0]pps$DMA1DRTYPE;
    wire pps$DMA1DRVALID;
    wire pps$DMA1RSTN;
    wire pps$DMA2ACLK;
    wire pps$DMA2DAREADY;
    wire [1:0]pps$DMA2DATYPE;
    wire pps$DMA2DAVALID;
    wire pps$DMA2DRLAST;
    wire pps$DMA2DRREADY;
    wire [1:0]pps$DMA2DRTYPE;
    wire pps$DMA2DRVALID;
    wire pps$DMA2RSTN;
    wire pps$DMA3ACLK;
    wire pps$DMA3DAREADY;
    wire [1:0]pps$DMA3DATYPE;
    wire pps$DMA3DAVALID;
    wire pps$DMA3DRLAST;
    wire pps$DMA3DRREADY;
    wire [1:0]pps$DMA3DRTYPE;
    wire pps$DMA3DRVALID;
    wire pps$DMA3RSTN;
    wire pps$EMIOCAN0PHYRX;
    wire pps$EMIOCAN0PHYTX;
    wire pps$EMIOCAN1PHYRX;
    wire pps$EMIOCAN1PHYTX;
    wire pps$EMIOENET0EXTINTIN;
    wire pps$EMIOENET0GMIICOL;
    wire pps$EMIOENET0GMIICRS;
    wire pps$EMIOENET0GMIIRXCLK;
    wire [7:0]pps$EMIOENET0GMIIRXD;
    wire pps$EMIOENET0GMIIRXDV;
    wire pps$EMIOENET0GMIIRXER;
    wire pps$EMIOENET0GMIITXCLK;
    wire [7:0]pps$EMIOENET0GMIITXD;
    wire pps$EMIOENET0GMIITXEN;
    wire pps$EMIOENET0GMIITXER;
    wire pps$EMIOENET0MDIOI;
    wire pps$EMIOENET0MDIOMDC;
    wire pps$EMIOENET0MDIOO;
    wire pps$EMIOENET0MDIOTN;
    wire pps$EMIOENET0PTPDELAYREQRX;
    wire pps$EMIOENET0PTPDELAYREQTX;
    wire pps$EMIOENET0PTPPDELAYREQRX;
    wire pps$EMIOENET0PTPPDELAYREQTX;
    wire pps$EMIOENET0PTPPDELAYRESPRX;
    wire pps$EMIOENET0PTPPDELAYRESPTX;
    wire pps$EMIOENET0PTPSYNCFRAMERX;
    wire pps$EMIOENET0PTPSYNCFRAMETX;
    wire pps$EMIOENET0SOFRX;
    wire pps$EMIOENET0SOFTX;
    wire pps$EMIOENET1EXTINTIN;
    wire pps$EMIOENET1GMIICOL;
    wire pps$EMIOENET1GMIICRS;
    wire pps$EMIOENET1GMIIRXCLK;
    wire [7:0]pps$EMIOENET1GMIIRXD;
    wire pps$EMIOENET1GMIIRXDV;
    wire pps$EMIOENET1GMIIRXER;
    wire pps$EMIOENET1GMIITXCLK;
    wire [7:0]pps$EMIOENET1GMIITXD;
    wire pps$EMIOENET1GMIITXEN;
    wire pps$EMIOENET1GMIITXER;
    wire pps$EMIOENET1MDIOI;
    wire pps$EMIOENET1MDIOMDC;
    wire pps$EMIOENET1MDIOO;
    wire pps$EMIOENET1MDIOTN;
    wire pps$EMIOENET1PTPDELAYREQRX;
    wire pps$EMIOENET1PTPDELAYREQTX;
    wire pps$EMIOENET1PTPPDELAYREQRX;
    wire pps$EMIOENET1PTPPDELAYREQTX;
    wire pps$EMIOENET1PTPPDELAYRESPRX;
    wire pps$EMIOENET1PTPPDELAYRESPTX;
    wire pps$EMIOENET1PTPSYNCFRAMERX;
    wire pps$EMIOENET1PTPSYNCFRAMETX;
    wire pps$EMIOENET1SOFRX;
    wire pps$EMIOENET1SOFTX;
    wire [63:0]pps$EMIOGPIOI;
    wire [63:0]pps$EMIOGPIOO;
    wire [63:0]pps$EMIOGPIOTN;
    wire pps$EMIOI2C0SCLI;
    wire pps$EMIOI2C0SCLO;
    wire pps$EMIOI2C0SCLTN;
    wire pps$EMIOI2C0SDAI;
    wire pps$EMIOI2C0SDAO;
    wire pps$EMIOI2C0SDATN;
    wire pps$EMIOI2C1SCLI;
    wire pps$EMIOI2C1SCLO;
    wire pps$EMIOI2C1SCLTN;
    wire pps$EMIOI2C1SDAI;
    wire pps$EMIOI2C1SDAO;
    wire pps$EMIOI2C1SDATN;
    wire pps$EMIOPJTAGTCK;
    wire pps$EMIOPJTAGTDI;
    wire pps$EMIOPJTAGTDO;
    wire pps$EMIOPJTAGTDTN;
    wire pps$EMIOPJTAGTMS;
    wire pps$EMIOSDIO0BUSPOW;
    wire [2:0]pps$EMIOSDIO0BUSVOLT;
    wire pps$EMIOSDIO0CDN;
    wire pps$EMIOSDIO0CLK;
    wire pps$EMIOSDIO0CLKFB;
    wire pps$EMIOSDIO0CMDI;
    wire pps$EMIOSDIO0CMDO;
    wire pps$EMIOSDIO0CMDTN;
    wire [3:0]pps$EMIOSDIO0DATAI;
    wire [3:0]pps$EMIOSDIO0DATAO;
    wire [3:0]pps$EMIOSDIO0DATATN;
    wire pps$EMIOSDIO0LED;
    wire pps$EMIOSDIO0WP;
    wire pps$EMIOSDIO1BUSPOW;
    wire [2:0]pps$EMIOSDIO1BUSVOLT;
    wire pps$EMIOSDIO1CDN;
    wire pps$EMIOSDIO1CLK;
    wire pps$EMIOSDIO1CLKFB;
    wire pps$EMIOSDIO1CMDI;
    wire pps$EMIOSDIO1CMDO;
    wire pps$EMIOSDIO1CMDTN;
    wire [3:0]pps$EMIOSDIO1DATAI;
    wire [3:0]pps$EMIOSDIO1DATAO;
    wire [3:0]pps$EMIOSDIO1DATATN;
    wire pps$EMIOSDIO1LED;
    wire pps$EMIOSDIO1WP;
    wire pps$EMIOSPI0MI;
    wire pps$EMIOSPI0MO;
    wire pps$EMIOSPI0MOTN;
    wire pps$EMIOSPI0SCLKI;
    wire pps$EMIOSPI0SCLKO;
    wire pps$EMIOSPI0SCLKTN;
    wire pps$EMIOSPI0SI;
    wire pps$EMIOSPI0SO;
    wire pps$EMIOSPI0SSIN;
    wire pps$EMIOSPI0SSNTN;
    wire [2:0]pps$EMIOSPI0SSON;
    wire pps$EMIOSPI0STN;
    wire pps$EMIOSPI1MI;
    wire pps$EMIOSPI1MO;
    wire pps$EMIOSPI1MOTN;
    wire pps$EMIOSPI1SCLKI;
    wire pps$EMIOSPI1SCLKO;
    wire pps$EMIOSPI1SCLKTN;
    wire pps$EMIOSPI1SI;
    wire pps$EMIOSPI1SO;
    wire pps$EMIOSPI1SSIN;
    wire pps$EMIOSPI1SSNTN;
    wire [2:0]pps$EMIOSPI1SSON;
    wire pps$EMIOSPI1STN;
    wire pps$EMIOSRAMINTIN;
    wire pps$EMIOTRACECLK;
    wire pps$EMIOTRACECTL;
    wire [31:0]pps$EMIOTRACEDATA;
    wire [2:0]pps$EMIOTTC0CLKI;
    wire [2:0]pps$EMIOTTC0WAVEO;
    wire [2:0]pps$EMIOTTC1CLKI;
    wire [2:0]pps$EMIOTTC1WAVEO;
    wire pps$EMIOUART0CTSN;
    wire pps$EMIOUART0DCDN;
    wire pps$EMIOUART0DSRN;
    wire pps$EMIOUART0DTRN;
    wire pps$EMIOUART0RIN;
    wire pps$EMIOUART0RTSN;
    wire pps$EMIOUART0RX;
    wire pps$EMIOUART0TX;
    wire pps$EMIOUART1CTSN;
    wire pps$EMIOUART1DCDN;
    wire pps$EMIOUART1DSRN;
    wire pps$EMIOUART1DTRN;
    wire pps$EMIOUART1RIN;
    wire pps$EMIOUART1RTSN;
    wire pps$EMIOUART1RX;
    wire pps$EMIOUART1TX;
    wire [1:0]pps$EMIOUSB0PORTINDCTL;
    wire pps$EMIOUSB0VBUSPWRFAULT;
    wire pps$EMIOUSB0VBUSPWRSELECT;
    wire [1:0]pps$EMIOUSB1PORTINDCTL;
    wire pps$EMIOUSB1VBUSPWRFAULT;
    wire pps$EMIOUSB1VBUSPWRSELECT;
    wire pps$EMIOWDTCLKI;
    wire pps$EMIOWDTRSTO;
    wire pps$EVENTEVENTI;
    wire pps$EVENTEVENTO;
    wire [1:0]pps$EVENTSTANDBYWFE;
    wire [1:0]pps$EVENTSTANDBYWFI;
    wire [3:0]pps$FCLKCLKTRIGN;
    wire [3:0]pps$FCLKRESETN;
    wire [3:0]pps$FTMDTRACEINATID;
    wire pps$FTMDTRACEINCLOCK;
    wire [31:0]pps$FTMDTRACEINDATA;
    wire pps$FTMDTRACEINVALID;
    wire [31:0]pps$FTMTF2PDEBUG;
    wire [3:0]pps$FTMTF2PTRIG;
    wire [3:0]pps$FTMTF2PTRIGACK;
    wire [31:0]pps$FTMTP2FDEBUG;
    wire [3:0]pps$FTMTP2FTRIG;
    wire [3:0]pps$FTMTP2FTRIGACK;
    wire [31:0]pps$MAXIGP1ARADDR;
    wire [1:0]pps$MAXIGP1ARBURST;
    wire [3:0]pps$MAXIGP1ARCACHE;
    wire pps$MAXIGP1ARESETN;
    wire [11:0]pps$MAXIGP1ARID;
    wire [3:0]pps$MAXIGP1ARLEN;
    wire [1:0]pps$MAXIGP1ARLOCK;
    wire [2:0]pps$MAXIGP1ARPROT;
    wire [3:0]pps$MAXIGP1ARQOS;
    wire pps$MAXIGP1ARREADY;
    wire [1:0]pps$MAXIGP1ARSIZE;
    wire pps$MAXIGP1ARVALID;
    wire [31:0]pps$MAXIGP1AWADDR;
    wire [1:0]pps$MAXIGP1AWBURST;
    wire [3:0]pps$MAXIGP1AWCACHE;
    wire [11:0]pps$MAXIGP1AWID;
    wire [3:0]pps$MAXIGP1AWLEN;
    wire [1:0]pps$MAXIGP1AWLOCK;
    wire [2:0]pps$MAXIGP1AWPROT;
    wire [3:0]pps$MAXIGP1AWQOS;
    wire pps$MAXIGP1AWREADY;
    wire [1:0]pps$MAXIGP1AWSIZE;
    wire pps$MAXIGP1AWVALID;
    wire [11:0]pps$MAXIGP1BID;
    wire pps$MAXIGP1BREADY;
    wire [1:0]pps$MAXIGP1BRESP;
    wire pps$MAXIGP1BVALID;
    wire [31:0]pps$MAXIGP1RDATA;
    wire [11:0]pps$MAXIGP1RID;
    wire pps$MAXIGP1RLAST;
    wire pps$MAXIGP1RREADY;
    wire [1:0]pps$MAXIGP1RRESP;
    wire pps$MAXIGP1RVALID;
    wire [31:0]pps$MAXIGP1WDATA;
    wire [11:0]pps$MAXIGP1WID;
    wire pps$MAXIGP1WLAST;
    wire pps$MAXIGP1WREADY;
    wire [3:0]pps$MAXIGP1WSTRB;
    wire pps$MAXIGP1WVALID;
    wire [31:0]pps$SAXIACPARADDR;
    wire [1:0]pps$SAXIACPARBURST;
    wire [3:0]pps$SAXIACPARCACHE;
    wire pps$SAXIACPARESETN;
    wire [2:0]pps$SAXIACPARID;
    wire [3:0]pps$SAXIACPARLEN;
    wire [1:0]pps$SAXIACPARLOCK;
    wire [2:0]pps$SAXIACPARPROT;
    wire [3:0]pps$SAXIACPARQOS;
    wire pps$SAXIACPARREADY;
    wire [1:0]pps$SAXIACPARSIZE;
    wire [4:0]pps$SAXIACPARUSER;
    wire pps$SAXIACPARVALID;
    wire [31:0]pps$SAXIACPAWADDR;
    wire [1:0]pps$SAXIACPAWBURST;
    wire [3:0]pps$SAXIACPAWCACHE;
    wire [2:0]pps$SAXIACPAWID;
    wire [3:0]pps$SAXIACPAWLEN;
    wire [1:0]pps$SAXIACPAWLOCK;
    wire [2:0]pps$SAXIACPAWPROT;
    wire [3:0]pps$SAXIACPAWQOS;
    wire pps$SAXIACPAWREADY;
    wire [1:0]pps$SAXIACPAWSIZE;
    wire [4:0]pps$SAXIACPAWUSER;
    wire pps$SAXIACPAWVALID;
    wire [2:0]pps$SAXIACPBID;
    wire pps$SAXIACPBREADY;
    wire [1:0]pps$SAXIACPBRESP;
    wire pps$SAXIACPBVALID;
    wire [63:0]pps$SAXIACPRDATA;
    wire [2:0]pps$SAXIACPRID;
    wire pps$SAXIACPRLAST;
    wire pps$SAXIACPRREADY;
    wire [1:0]pps$SAXIACPRRESP;
    wire pps$SAXIACPRVALID;
    wire [63:0]pps$SAXIACPWDATA;
    wire [2:0]pps$SAXIACPWID;
    wire pps$SAXIACPWLAST;
    wire pps$SAXIACPWREADY;
    wire [7:0]pps$SAXIACPWSTRB;
    wire pps$SAXIACPWVALID;
    wire [31:0]pps$SAXIGP0ARADDR;
    wire [1:0]pps$SAXIGP0ARBURST;
    wire [3:0]pps$SAXIGP0ARCACHE;
    wire pps$SAXIGP0ARESETN;
    wire [5:0]pps$SAXIGP0ARID;
    wire [3:0]pps$SAXIGP0ARLEN;
    wire [1:0]pps$SAXIGP0ARLOCK;
    wire [2:0]pps$SAXIGP0ARPROT;
    wire [3:0]pps$SAXIGP0ARQOS;
    wire pps$SAXIGP0ARREADY;
    wire [1:0]pps$SAXIGP0ARSIZE;
    wire pps$SAXIGP0ARVALID;
    wire [31:0]pps$SAXIGP0AWADDR;
    wire [1:0]pps$SAXIGP0AWBURST;
    wire [3:0]pps$SAXIGP0AWCACHE;
    wire [5:0]pps$SAXIGP0AWID;
    wire [3:0]pps$SAXIGP0AWLEN;
    wire [1:0]pps$SAXIGP0AWLOCK;
    wire [2:0]pps$SAXIGP0AWPROT;
    wire [3:0]pps$SAXIGP0AWQOS;
    wire pps$SAXIGP0AWREADY;
    wire [1:0]pps$SAXIGP0AWSIZE;
    wire pps$SAXIGP0AWVALID;
    wire [5:0]pps$SAXIGP0BID;
    wire pps$SAXIGP0BREADY;
    wire [1:0]pps$SAXIGP0BRESP;
    wire pps$SAXIGP0BVALID;
    wire [31:0]pps$SAXIGP0RDATA;
    wire [5:0]pps$SAXIGP0RID;
    wire pps$SAXIGP0RLAST;
    wire pps$SAXIGP0RREADY;
    wire [1:0]pps$SAXIGP0RRESP;
    wire pps$SAXIGP0RVALID;
    wire [31:0]pps$SAXIGP0WDATA;
    wire [5:0]pps$SAXIGP0WID;
    wire pps$SAXIGP0WLAST;
    wire pps$SAXIGP0WREADY;
    wire [3:0]pps$SAXIGP0WSTRB;
    wire pps$SAXIGP0WVALID;
    wire [31:0]pps$SAXIGP1ARADDR;
    wire [1:0]pps$SAXIGP1ARBURST;
    wire [3:0]pps$SAXIGP1ARCACHE;
    wire pps$SAXIGP1ARESETN;
    wire [5:0]pps$SAXIGP1ARID;
    wire [3:0]pps$SAXIGP1ARLEN;
    wire [1:0]pps$SAXIGP1ARLOCK;
    wire [2:0]pps$SAXIGP1ARPROT;
    wire [3:0]pps$SAXIGP1ARQOS;
    wire pps$SAXIGP1ARREADY;
    wire [1:0]pps$SAXIGP1ARSIZE;
    wire pps$SAXIGP1ARVALID;
    wire [31:0]pps$SAXIGP1AWADDR;
    wire [1:0]pps$SAXIGP1AWBURST;
    wire [3:0]pps$SAXIGP1AWCACHE;
    wire [5:0]pps$SAXIGP1AWID;
    wire [3:0]pps$SAXIGP1AWLEN;
    wire [1:0]pps$SAXIGP1AWLOCK;
    wire [2:0]pps$SAXIGP1AWPROT;
    wire [3:0]pps$SAXIGP1AWQOS;
    wire pps$SAXIGP1AWREADY;
    wire [1:0]pps$SAXIGP1AWSIZE;
    wire pps$SAXIGP1AWVALID;
    wire [5:0]pps$SAXIGP1BID;
    wire pps$SAXIGP1BREADY;
    wire [1:0]pps$SAXIGP1BRESP;
    wire pps$SAXIGP1BVALID;
    wire [31:0]pps$SAXIGP1RDATA;
    wire [5:0]pps$SAXIGP1RID;
    wire pps$SAXIGP1RLAST;
    wire pps$SAXIGP1RREADY;
    wire [1:0]pps$SAXIGP1RRESP;
    wire pps$SAXIGP1RVALID;
    wire [31:0]pps$SAXIGP1WDATA;
    wire [5:0]pps$SAXIGP1WID;
    wire pps$SAXIGP1WLAST;
    wire pps$SAXIGP1WREADY;
    wire [3:0]pps$SAXIGP1WSTRB;
    wire pps$SAXIGP1WVALID;
    wire [31:0]pps$SAXIHP0ARADDR;
    wire [1:0]pps$SAXIHP0ARBURST;
    wire [3:0]pps$SAXIHP0ARCACHE;
    wire pps$SAXIHP0ARESETN;
    wire [5:0]pps$SAXIHP0ARID;
    wire [3:0]pps$SAXIHP0ARLEN;
    wire [1:0]pps$SAXIHP0ARLOCK;
    wire [2:0]pps$SAXIHP0ARPROT;
    wire [3:0]pps$SAXIHP0ARQOS;
    wire pps$SAXIHP0ARREADY;
    wire [1:0]pps$SAXIHP0ARSIZE;
    wire pps$SAXIHP0ARVALID;
    wire [31:0]pps$SAXIHP0AWADDR;
    wire [1:0]pps$SAXIHP0AWBURST;
    wire [3:0]pps$SAXIHP0AWCACHE;
    wire [5:0]pps$SAXIHP0AWID;
    wire [3:0]pps$SAXIHP0AWLEN;
    wire [1:0]pps$SAXIHP0AWLOCK;
    wire [2:0]pps$SAXIHP0AWPROT;
    wire [3:0]pps$SAXIHP0AWQOS;
    wire pps$SAXIHP0AWREADY;
    wire [1:0]pps$SAXIHP0AWSIZE;
    wire pps$SAXIHP0AWVALID;
    wire [5:0]pps$SAXIHP0BID;
    wire pps$SAXIHP0BREADY;
    wire [1:0]pps$SAXIHP0BRESP;
    wire pps$SAXIHP0BVALID;
    wire [2:0]pps$SAXIHP0RACOUNT;
    wire [7:0]pps$SAXIHP0RCOUNT;
    wire [63:0]pps$SAXIHP0RDATA;
    wire pps$SAXIHP0RDISSUECAP1EN;
    wire [5:0]pps$SAXIHP0RID;
    wire pps$SAXIHP0RLAST;
    wire pps$SAXIHP0RREADY;
    wire [1:0]pps$SAXIHP0RRESP;
    wire pps$SAXIHP0RVALID;
    wire [5:0]pps$SAXIHP0WACOUNT;
    wire [7:0]pps$SAXIHP0WCOUNT;
    wire [63:0]pps$SAXIHP0WDATA;
    wire [5:0]pps$SAXIHP0WID;
    wire pps$SAXIHP0WLAST;
    wire pps$SAXIHP0WREADY;
    wire pps$SAXIHP0WRISSUECAP1EN;
    wire [7:0]pps$SAXIHP0WSTRB;
    wire pps$SAXIHP0WVALID;
    wire [31:0]pps$SAXIHP1ARADDR;
    wire [1:0]pps$SAXIHP1ARBURST;
    wire [3:0]pps$SAXIHP1ARCACHE;
    wire pps$SAXIHP1ARESETN;
    wire [5:0]pps$SAXIHP1ARID;
    wire [3:0]pps$SAXIHP1ARLEN;
    wire [1:0]pps$SAXIHP1ARLOCK;
    wire [2:0]pps$SAXIHP1ARPROT;
    wire [3:0]pps$SAXIHP1ARQOS;
    wire pps$SAXIHP1ARREADY;
    wire [1:0]pps$SAXIHP1ARSIZE;
    wire pps$SAXIHP1ARVALID;
    wire [31:0]pps$SAXIHP1AWADDR;
    wire [1:0]pps$SAXIHP1AWBURST;
    wire [3:0]pps$SAXIHP1AWCACHE;
    wire [5:0]pps$SAXIHP1AWID;
    wire [3:0]pps$SAXIHP1AWLEN;
    wire [1:0]pps$SAXIHP1AWLOCK;
    wire [2:0]pps$SAXIHP1AWPROT;
    wire [3:0]pps$SAXIHP1AWQOS;
    wire pps$SAXIHP1AWREADY;
    wire [1:0]pps$SAXIHP1AWSIZE;
    wire pps$SAXIHP1AWVALID;
    wire [5:0]pps$SAXIHP1BID;
    wire pps$SAXIHP1BREADY;
    wire [1:0]pps$SAXIHP1BRESP;
    wire pps$SAXIHP1BVALID;
    wire [2:0]pps$SAXIHP1RACOUNT;
    wire [7:0]pps$SAXIHP1RCOUNT;
    wire [63:0]pps$SAXIHP1RDATA;
    wire pps$SAXIHP1RDISSUECAP1EN;
    wire [5:0]pps$SAXIHP1RID;
    wire pps$SAXIHP1RLAST;
    wire pps$SAXIHP1RREADY;
    wire [1:0]pps$SAXIHP1RRESP;
    wire pps$SAXIHP1RVALID;
    wire [5:0]pps$SAXIHP1WACOUNT;
    wire [7:0]pps$SAXIHP1WCOUNT;
    wire [63:0]pps$SAXIHP1WDATA;
    wire [5:0]pps$SAXIHP1WID;
    wire pps$SAXIHP1WLAST;
    wire pps$SAXIHP1WREADY;
    wire pps$SAXIHP1WRISSUECAP1EN;
    wire [7:0]pps$SAXIHP1WSTRB;
    wire pps$SAXIHP1WVALID;
    wire [31:0]pps$SAXIHP2ARADDR;
    wire [1:0]pps$SAXIHP2ARBURST;
    wire [3:0]pps$SAXIHP2ARCACHE;
    wire pps$SAXIHP2ARESETN;
    wire [5:0]pps$SAXIHP2ARID;
    wire [3:0]pps$SAXIHP2ARLEN;
    wire [1:0]pps$SAXIHP2ARLOCK;
    wire [2:0]pps$SAXIHP2ARPROT;
    wire [3:0]pps$SAXIHP2ARQOS;
    wire pps$SAXIHP2ARREADY;
    wire [1:0]pps$SAXIHP2ARSIZE;
    wire pps$SAXIHP2ARVALID;
    wire [31:0]pps$SAXIHP2AWADDR;
    wire [1:0]pps$SAXIHP2AWBURST;
    wire [3:0]pps$SAXIHP2AWCACHE;
    wire [5:0]pps$SAXIHP2AWID;
    wire [3:0]pps$SAXIHP2AWLEN;
    wire [1:0]pps$SAXIHP2AWLOCK;
    wire [2:0]pps$SAXIHP2AWPROT;
    wire [3:0]pps$SAXIHP2AWQOS;
    wire pps$SAXIHP2AWREADY;
    wire [1:0]pps$SAXIHP2AWSIZE;
    wire pps$SAXIHP2AWVALID;
    wire [5:0]pps$SAXIHP2BID;
    wire pps$SAXIHP2BREADY;
    wire [1:0]pps$SAXIHP2BRESP;
    wire pps$SAXIHP2BVALID;
    wire [2:0]pps$SAXIHP2RACOUNT;
    wire [7:0]pps$SAXIHP2RCOUNT;
    wire [63:0]pps$SAXIHP2RDATA;
    wire pps$SAXIHP2RDISSUECAP1EN;
    wire [5:0]pps$SAXIHP2RID;
    wire pps$SAXIHP2RLAST;
    wire pps$SAXIHP2RREADY;
    wire [1:0]pps$SAXIHP2RRESP;
    wire pps$SAXIHP2RVALID;
    wire [5:0]pps$SAXIHP2WACOUNT;
    wire [7:0]pps$SAXIHP2WCOUNT;
    wire [63:0]pps$SAXIHP2WDATA;
    wire [5:0]pps$SAXIHP2WID;
    wire pps$SAXIHP2WLAST;
    wire pps$SAXIHP2WREADY;
    wire pps$SAXIHP2WRISSUECAP1EN;
    wire [7:0]pps$SAXIHP2WSTRB;
    wire pps$SAXIHP2WVALID;
    wire [31:0]pps$SAXIHP3ARADDR;
    wire [1:0]pps$SAXIHP3ARBURST;
    wire [3:0]pps$SAXIHP3ARCACHE;
    wire pps$SAXIHP3ARESETN;
    wire [5:0]pps$SAXIHP3ARID;
    wire [3:0]pps$SAXIHP3ARLEN;
    wire [1:0]pps$SAXIHP3ARLOCK;
    wire [2:0]pps$SAXIHP3ARPROT;
    wire [3:0]pps$SAXIHP3ARQOS;
    wire pps$SAXIHP3ARREADY;
    wire [1:0]pps$SAXIHP3ARSIZE;
    wire pps$SAXIHP3ARVALID;
    wire [31:0]pps$SAXIHP3AWADDR;
    wire [1:0]pps$SAXIHP3AWBURST;
    wire [3:0]pps$SAXIHP3AWCACHE;
    wire [5:0]pps$SAXIHP3AWID;
    wire [3:0]pps$SAXIHP3AWLEN;
    wire [1:0]pps$SAXIHP3AWLOCK;
    wire [2:0]pps$SAXIHP3AWPROT;
    wire [3:0]pps$SAXIHP3AWQOS;
    wire pps$SAXIHP3AWREADY;
    wire [1:0]pps$SAXIHP3AWSIZE;
    wire pps$SAXIHP3AWVALID;
    wire [5:0]pps$SAXIHP3BID;
    wire pps$SAXIHP3BREADY;
    wire [1:0]pps$SAXIHP3BRESP;
    wire pps$SAXIHP3BVALID;
    wire [2:0]pps$SAXIHP3RACOUNT;
    wire [7:0]pps$SAXIHP3RCOUNT;
    wire [63:0]pps$SAXIHP3RDATA;
    wire pps$SAXIHP3RDISSUECAP1EN;
    wire [5:0]pps$SAXIHP3RID;
    wire pps$SAXIHP3RLAST;
    wire pps$SAXIHP3RREADY;
    wire [1:0]pps$SAXIHP3RRESP;
    wire pps$SAXIHP3RVALID;
    wire [5:0]pps$SAXIHP3WACOUNT;
    wire [7:0]pps$SAXIHP3WCOUNT;
    wire [63:0]pps$SAXIHP3WDATA;
    wire [5:0]pps$SAXIHP3WID;
    wire pps$SAXIHP3WLAST;
    wire pps$SAXIHP3WREADY;
    wire pps$SAXIHP3WRISSUECAP1EN;
    wire [7:0]pps$SAXIHP3WSTRB;
    wire pps$SAXIHP3WVALID;
    assign init__ENA = 1;
    PS7 pps (
        .DDRA(DDRA),
        .DDRARB(DDRARB),
        .DDRBA(DDRBA),
        .DDRCASB(DDRCASB),
        .DDRCKE(DDRCKE),
        .DDRCKN(DDRCKN),
        .DDRCKP(DDRCKP),
        .DDRCSB(DDRCSB),
        .DDRDM(DDRDM),
        .DDRDQ(DDRDQ),
        .DDRDQSN(DDRDQSN),
        .DDRDQSP(DDRDQSP),
        .DDRDRSTB(DDRDRSTB),
        .DDRODT(DDRODT),
        .DDRRASB(DDRRASB),
        .DDRVRN(DDRVRN),
        .DDRVRP(DDRVRP),
        .DDRWEB(DDRWEB),
        .DMA0ACLK(pps$DMA0ACLK),
        .DMA0DAREADY(pps$DMA0DAREADY),
        .DMA0DATYPE(pps$DMA0DATYPE),
        .DMA0DAVALID(pps$DMA0DAVALID),
        .DMA0DRLAST(pps$DMA0DRLAST),
        .DMA0DRREADY(pps$DMA0DRREADY),
        .DMA0DRTYPE(pps$DMA0DRTYPE),
        .DMA0DRVALID(pps$DMA0DRVALID),
        .DMA0RSTN(pps$DMA0RSTN),
        .DMA1ACLK(pps$DMA1ACLK),
        .DMA1DAREADY(pps$DMA1DAREADY),
        .DMA1DATYPE(pps$DMA1DATYPE),
        .DMA1DAVALID(pps$DMA1DAVALID),
        .DMA1DRLAST(pps$DMA1DRLAST),
        .DMA1DRREADY(pps$DMA1DRREADY),
        .DMA1DRTYPE(pps$DMA1DRTYPE),
        .DMA1DRVALID(pps$DMA1DRVALID),
        .DMA1RSTN(pps$DMA1RSTN),
        .DMA2ACLK(pps$DMA2ACLK),
        .DMA2DAREADY(pps$DMA2DAREADY),
        .DMA2DATYPE(pps$DMA2DATYPE),
        .DMA2DAVALID(pps$DMA2DAVALID),
        .DMA2DRLAST(pps$DMA2DRLAST),
        .DMA2DRREADY(pps$DMA2DRREADY),
        .DMA2DRTYPE(pps$DMA2DRTYPE),
        .DMA2DRVALID(pps$DMA2DRVALID),
        .DMA2RSTN(pps$DMA2RSTN),
        .DMA3ACLK(pps$DMA3ACLK),
        .DMA3DAREADY(pps$DMA3DAREADY),
        .DMA3DATYPE(pps$DMA3DATYPE),
        .DMA3DAVALID(pps$DMA3DAVALID),
        .DMA3DRLAST(pps$DMA3DRLAST),
        .DMA3DRREADY(pps$DMA3DRREADY),
        .DMA3DRTYPE(pps$DMA3DRTYPE),
        .DMA3DRVALID(pps$DMA3DRVALID),
        .DMA3RSTN(pps$DMA3RSTN),
        .EMIOCAN0PHYRX(pps$EMIOCAN0PHYRX),
        .EMIOCAN0PHYTX(pps$EMIOCAN0PHYTX),
        .EMIOCAN1PHYRX(pps$EMIOCAN1PHYRX),
        .EMIOCAN1PHYTX(pps$EMIOCAN1PHYTX),
        .EMIOENET0EXTINTIN(pps$EMIOENET0EXTINTIN),
        .EMIOENET0GMIICOL(pps$EMIOENET0GMIICOL),
        .EMIOENET0GMIICRS(pps$EMIOENET0GMIICRS),
        .EMIOENET0GMIIRXCLK(pps$EMIOENET0GMIIRXCLK),
        .EMIOENET0GMIIRXD(pps$EMIOENET0GMIIRXD),
        .EMIOENET0GMIIRXDV(pps$EMIOENET0GMIIRXDV),
        .EMIOENET0GMIIRXER(pps$EMIOENET0GMIIRXER),
        .EMIOENET0GMIITXCLK(pps$EMIOENET0GMIITXCLK),
        .EMIOENET0GMIITXD(pps$EMIOENET0GMIITXD),
        .EMIOENET0GMIITXEN(pps$EMIOENET0GMIITXEN),
        .EMIOENET0GMIITXER(pps$EMIOENET0GMIITXER),
        .EMIOENET0MDIOI(pps$EMIOENET0MDIOI),
        .EMIOENET0MDIOMDC(pps$EMIOENET0MDIOMDC),
        .EMIOENET0MDIOO(pps$EMIOENET0MDIOO),
        .EMIOENET0MDIOTN(pps$EMIOENET0MDIOTN),
        .EMIOENET0PTPDELAYREQRX(pps$EMIOENET0PTPDELAYREQRX),
        .EMIOENET0PTPDELAYREQTX(pps$EMIOENET0PTPDELAYREQTX),
        .EMIOENET0PTPPDELAYREQRX(pps$EMIOENET0PTPPDELAYREQRX),
        .EMIOENET0PTPPDELAYREQTX(pps$EMIOENET0PTPPDELAYREQTX),
        .EMIOENET0PTPPDELAYRESPRX(pps$EMIOENET0PTPPDELAYRESPRX),
        .EMIOENET0PTPPDELAYRESPTX(pps$EMIOENET0PTPPDELAYRESPTX),
        .EMIOENET0PTPSYNCFRAMERX(pps$EMIOENET0PTPSYNCFRAMERX),
        .EMIOENET0PTPSYNCFRAMETX(pps$EMIOENET0PTPSYNCFRAMETX),
        .EMIOENET0SOFRX(pps$EMIOENET0SOFRX),
        .EMIOENET0SOFTX(pps$EMIOENET0SOFTX),
        .EMIOENET1EXTINTIN(pps$EMIOENET1EXTINTIN),
        .EMIOENET1GMIICOL(pps$EMIOENET1GMIICOL),
        .EMIOENET1GMIICRS(pps$EMIOENET1GMIICRS),
        .EMIOENET1GMIIRXCLK(pps$EMIOENET1GMIIRXCLK),
        .EMIOENET1GMIIRXD(pps$EMIOENET1GMIIRXD),
        .EMIOENET1GMIIRXDV(pps$EMIOENET1GMIIRXDV),
        .EMIOENET1GMIIRXER(pps$EMIOENET1GMIIRXER),
        .EMIOENET1GMIITXCLK(pps$EMIOENET1GMIITXCLK),
        .EMIOENET1GMIITXD(pps$EMIOENET1GMIITXD),
        .EMIOENET1GMIITXEN(pps$EMIOENET1GMIITXEN),
        .EMIOENET1GMIITXER(pps$EMIOENET1GMIITXER),
        .EMIOENET1MDIOI(pps$EMIOENET1MDIOI),
        .EMIOENET1MDIOMDC(pps$EMIOENET1MDIOMDC),
        .EMIOENET1MDIOO(pps$EMIOENET1MDIOO),
        .EMIOENET1MDIOTN(pps$EMIOENET1MDIOTN),
        .EMIOENET1PTPDELAYREQRX(pps$EMIOENET1PTPDELAYREQRX),
        .EMIOENET1PTPDELAYREQTX(pps$EMIOENET1PTPDELAYREQTX),
        .EMIOENET1PTPPDELAYREQRX(pps$EMIOENET1PTPPDELAYREQRX),
        .EMIOENET1PTPPDELAYREQTX(pps$EMIOENET1PTPPDELAYREQTX),
        .EMIOENET1PTPPDELAYRESPRX(pps$EMIOENET1PTPPDELAYRESPRX),
        .EMIOENET1PTPPDELAYRESPTX(pps$EMIOENET1PTPPDELAYRESPTX),
        .EMIOENET1PTPSYNCFRAMERX(pps$EMIOENET1PTPSYNCFRAMERX),
        .EMIOENET1PTPSYNCFRAMETX(pps$EMIOENET1PTPSYNCFRAMETX),
        .EMIOENET1SOFRX(pps$EMIOENET1SOFRX),
        .EMIOENET1SOFTX(pps$EMIOENET1SOFTX),
        .EMIOGPIOI(pps$EMIOGPIOI),
        .EMIOGPIOO(pps$EMIOGPIOO),
        .EMIOGPIOTN(pps$EMIOGPIOTN),
        .EMIOI2C0SCLI(pps$EMIOI2C0SCLI),
        .EMIOI2C0SCLO(pps$EMIOI2C0SCLO),
        .EMIOI2C0SCLTN(pps$EMIOI2C0SCLTN),
        .EMIOI2C0SDAI(pps$EMIOI2C0SDAI),
        .EMIOI2C0SDAO(pps$EMIOI2C0SDAO),
        .EMIOI2C0SDATN(pps$EMIOI2C0SDATN),
        .EMIOI2C1SCLI(pps$EMIOI2C1SCLI),
        .EMIOI2C1SCLO(pps$EMIOI2C1SCLO),
        .EMIOI2C1SCLTN(pps$EMIOI2C1SCLTN),
        .EMIOI2C1SDAI(pps$EMIOI2C1SDAI),
        .EMIOI2C1SDAO(pps$EMIOI2C1SDAO),
        .EMIOI2C1SDATN(pps$EMIOI2C1SDATN),
        .EMIOPJTAGTCK(pps$EMIOPJTAGTCK),
        .EMIOPJTAGTDI(pps$EMIOPJTAGTDI),
        .EMIOPJTAGTDO(pps$EMIOPJTAGTDO),
        .EMIOPJTAGTDTN(pps$EMIOPJTAGTDTN),
        .EMIOPJTAGTMS(pps$EMIOPJTAGTMS),
        .EMIOSDIO0BUSPOW(pps$EMIOSDIO0BUSPOW),
        .EMIOSDIO0BUSVOLT(pps$EMIOSDIO0BUSVOLT),
        .EMIOSDIO0CDN(pps$EMIOSDIO0CDN),
        .EMIOSDIO0CLK(pps$EMIOSDIO0CLK),
        .EMIOSDIO0CLKFB(pps$EMIOSDIO0CLKFB),
        .EMIOSDIO0CMDI(pps$EMIOSDIO0CMDI),
        .EMIOSDIO0CMDO(pps$EMIOSDIO0CMDO),
        .EMIOSDIO0CMDTN(pps$EMIOSDIO0CMDTN),
        .EMIOSDIO0DATAI(pps$EMIOSDIO0DATAI),
        .EMIOSDIO0DATAO(pps$EMIOSDIO0DATAO),
        .EMIOSDIO0DATATN(pps$EMIOSDIO0DATATN),
        .EMIOSDIO0LED(pps$EMIOSDIO0LED),
        .EMIOSDIO0WP(pps$EMIOSDIO0WP),
        .EMIOSDIO1BUSPOW(pps$EMIOSDIO1BUSPOW),
        .EMIOSDIO1BUSVOLT(pps$EMIOSDIO1BUSVOLT),
        .EMIOSDIO1CDN(pps$EMIOSDIO1CDN),
        .EMIOSDIO1CLK(pps$EMIOSDIO1CLK),
        .EMIOSDIO1CLKFB(pps$EMIOSDIO1CLKFB),
        .EMIOSDIO1CMDI(pps$EMIOSDIO1CMDI),
        .EMIOSDIO1CMDO(pps$EMIOSDIO1CMDO),
        .EMIOSDIO1CMDTN(pps$EMIOSDIO1CMDTN),
        .EMIOSDIO1DATAI(pps$EMIOSDIO1DATAI),
        .EMIOSDIO1DATAO(pps$EMIOSDIO1DATAO),
        .EMIOSDIO1DATATN(pps$EMIOSDIO1DATATN),
        .EMIOSDIO1LED(pps$EMIOSDIO1LED),
        .EMIOSDIO1WP(pps$EMIOSDIO1WP),
        .EMIOSPI0MI(pps$EMIOSPI0MI),
        .EMIOSPI0MO(pps$EMIOSPI0MO),
        .EMIOSPI0MOTN(pps$EMIOSPI0MOTN),
        .EMIOSPI0SCLKI(pps$EMIOSPI0SCLKI),
        .EMIOSPI0SCLKO(pps$EMIOSPI0SCLKO),
        .EMIOSPI0SCLKTN(pps$EMIOSPI0SCLKTN),
        .EMIOSPI0SI(pps$EMIOSPI0SI),
        .EMIOSPI0SO(pps$EMIOSPI0SO),
        .EMIOSPI0SSIN(pps$EMIOSPI0SSIN),
        .EMIOSPI0SSNTN(pps$EMIOSPI0SSNTN),
        .EMIOSPI0SSON(pps$EMIOSPI0SSON),
        .EMIOSPI0STN(pps$EMIOSPI0STN),
        .EMIOSPI1MI(pps$EMIOSPI1MI),
        .EMIOSPI1MO(pps$EMIOSPI1MO),
        .EMIOSPI1MOTN(pps$EMIOSPI1MOTN),
        .EMIOSPI1SCLKI(pps$EMIOSPI1SCLKI),
        .EMIOSPI1SCLKO(pps$EMIOSPI1SCLKO),
        .EMIOSPI1SCLKTN(pps$EMIOSPI1SCLKTN),
        .EMIOSPI1SI(pps$EMIOSPI1SI),
        .EMIOSPI1SO(pps$EMIOSPI1SO),
        .EMIOSPI1SSIN(pps$EMIOSPI1SSIN),
        .EMIOSPI1SSNTN(pps$EMIOSPI1SSNTN),
        .EMIOSPI1SSON(pps$EMIOSPI1SSON),
        .EMIOSPI1STN(pps$EMIOSPI1STN),
        .EMIOSRAMINTIN(pps$EMIOSRAMINTIN),
        .EMIOTRACECLK(pps$EMIOTRACECLK),
        .EMIOTRACECTL(pps$EMIOTRACECTL),
        .EMIOTRACEDATA(pps$EMIOTRACEDATA),
        .EMIOTTC0CLKI(pps$EMIOTTC0CLKI),
        .EMIOTTC0WAVEO(pps$EMIOTTC0WAVEO),
        .EMIOTTC1CLKI(pps$EMIOTTC1CLKI),
        .EMIOTTC1WAVEO(pps$EMIOTTC1WAVEO),
        .EMIOUART0CTSN(pps$EMIOUART0CTSN),
        .EMIOUART0DCDN(pps$EMIOUART0DCDN),
        .EMIOUART0DSRN(pps$EMIOUART0DSRN),
        .EMIOUART0DTRN(pps$EMIOUART0DTRN),
        .EMIOUART0RIN(pps$EMIOUART0RIN),
        .EMIOUART0RTSN(pps$EMIOUART0RTSN),
        .EMIOUART0RX(pps$EMIOUART0RX),
        .EMIOUART0TX(pps$EMIOUART0TX),
        .EMIOUART1CTSN(pps$EMIOUART1CTSN),
        .EMIOUART1DCDN(pps$EMIOUART1DCDN),
        .EMIOUART1DSRN(pps$EMIOUART1DSRN),
        .EMIOUART1DTRN(pps$EMIOUART1DTRN),
        .EMIOUART1RIN(pps$EMIOUART1RIN),
        .EMIOUART1RTSN(pps$EMIOUART1RTSN),
        .EMIOUART1RX(pps$EMIOUART1RX),
        .EMIOUART1TX(pps$EMIOUART1TX),
        .EMIOUSB0PORTINDCTL(pps$EMIOUSB0PORTINDCTL),
        .EMIOUSB0VBUSPWRFAULT(pps$EMIOUSB0VBUSPWRFAULT),
        .EMIOUSB0VBUSPWRSELECT(pps$EMIOUSB0VBUSPWRSELECT),
        .EMIOUSB1PORTINDCTL(pps$EMIOUSB1PORTINDCTL),
        .EMIOUSB1VBUSPWRFAULT(pps$EMIOUSB1VBUSPWRFAULT),
        .EMIOUSB1VBUSPWRSELECT(pps$EMIOUSB1VBUSPWRSELECT),
        .EMIOWDTCLKI(pps$EMIOWDTCLKI),
        .EMIOWDTRSTO(pps$EMIOWDTRSTO),
        .EVENTEVENTI(pps$EVENTEVENTI),
        .EVENTEVENTO(pps$EVENTEVENTO),
        .EVENTSTANDBYWFE(pps$EVENTSTANDBYWFE),
        .EVENTSTANDBYWFI(pps$EVENTSTANDBYWFI),
        .FCLKCLK(FCLKCLK),
        .FCLKCLKTRIGN(pps$FCLKCLKTRIGN),
        .FCLKRESETN(pps$FCLKRESETN),
        .FPGAIDLEN(1'd1),
        .FTMDTRACEINATID(pps$FTMDTRACEINATID),
        .FTMDTRACEINCLOCK(pps$FTMDTRACEINCLOCK),
        .FTMDTRACEINDATA(pps$FTMDTRACEINDATA),
        .FTMDTRACEINVALID(pps$FTMDTRACEINVALID),
        .FTMTF2PDEBUG(pps$FTMTF2PDEBUG),
        .FTMTF2PTRIG(pps$FTMTF2PTRIG),
        .FTMTF2PTRIGACK(pps$FTMTF2PTRIGACK),
        .FTMTP2FDEBUG(pps$FTMTP2FDEBUG),
        .FTMTP2FTRIG(pps$FTMTP2FTRIG),
        .FTMTP2FTRIGACK(pps$FTMTP2FTRIGACK),
        .IRQF2P(IRQF2P),
        .IRQP2F(IRQP2F),
        .MAXIGP0ACLK(MAXIGP0ACLK),
        .MAXIGP0ARADDR(MAXIGP0ARADDR),
        .MAXIGP0ARBURST(MAXIGP0ARBURST),
        .MAXIGP0ARCACHE(MAXIGP0ARCACHE),
        .MAXIGP0ARESETN(MAXIGP0ARESETN),
        .MAXIGP0ARID(MAXIGP0ARID),
        .MAXIGP0ARLEN(MAXIGP0ARLEN),
        .MAXIGP0ARLOCK(MAXIGP0ARLOCK),
        .MAXIGP0ARPROT(MAXIGP0ARPROT),
        .MAXIGP0ARQOS(MAXIGP0ARQOS),
        .MAXIGP0ARREADY(MAXIGP0ARREADY),
        .MAXIGP0ARSIZE(MAXIGP0ARSIZE),
        .MAXIGP0ARVALID(MAXIGP0ARVALID),
        .MAXIGP0AWADDR(MAXIGP0AWADDR),
        .MAXIGP0AWBURST(MAXIGP0AWBURST),
        .MAXIGP0AWCACHE(MAXIGP0AWCACHE),
        .MAXIGP0AWID(MAXIGP0AWID),
        .MAXIGP0AWLEN(MAXIGP0AWLEN),
        .MAXIGP0AWLOCK(MAXIGP0AWLOCK),
        .MAXIGP0AWPROT(MAXIGP0AWPROT),
        .MAXIGP0AWQOS(MAXIGP0AWQOS),
        .MAXIGP0AWREADY(MAXIGP0AWREADY),
        .MAXIGP0AWSIZE(MAXIGP0AWSIZE),
        .MAXIGP0AWVALID(MAXIGP0AWVALID),
        .MAXIGP0BID(MAXIGP0BID),
        .MAXIGP0BREADY(MAXIGP0BREADY),
        .MAXIGP0BRESP(MAXIGP0BRESP),
        .MAXIGP0BVALID(MAXIGP0BVALID),
        .MAXIGP0RDATA(MAXIGP0RDATA),
        .MAXIGP0RID(MAXIGP0RID),
        .MAXIGP0RLAST(MAXIGP0RLAST),
        .MAXIGP0RREADY(MAXIGP0RREADY),
        .MAXIGP0RRESP(MAXIGP0RRESP),
        .MAXIGP0RVALID(MAXIGP0RVALID),
        .MAXIGP0WDATA(MAXIGP0WDATA),
        .MAXIGP0WID(MAXIGP0WID),
        .MAXIGP0WLAST(MAXIGP0WLAST),
        .MAXIGP0WREADY(MAXIGP0WREADY),
        .MAXIGP0WSTRB(MAXIGP0WSTRB),
        .MAXIGP0WVALID(MAXIGP0WVALID),
        .MAXIGP1ACLK(CLK),
        .MAXIGP1ARADDR(pps$MAXIGP1ARADDR),
        .MAXIGP1ARBURST(pps$MAXIGP1ARBURST),
        .MAXIGP1ARCACHE(pps$MAXIGP1ARCACHE),
        .MAXIGP1ARESETN(pps$MAXIGP1ARESETN),
        .MAXIGP1ARID(pps$MAXIGP1ARID),
        .MAXIGP1ARLEN(pps$MAXIGP1ARLEN),
        .MAXIGP1ARLOCK(pps$MAXIGP1ARLOCK),
        .MAXIGP1ARPROT(pps$MAXIGP1ARPROT),
        .MAXIGP1ARQOS(pps$MAXIGP1ARQOS),
        .MAXIGP1ARREADY(pps$MAXIGP1ARREADY),
        .MAXIGP1ARSIZE(pps$MAXIGP1ARSIZE),
        .MAXIGP1ARVALID(pps$MAXIGP1ARVALID),
        .MAXIGP1AWADDR(pps$MAXIGP1AWADDR),
        .MAXIGP1AWBURST(pps$MAXIGP1AWBURST),
        .MAXIGP1AWCACHE(pps$MAXIGP1AWCACHE),
        .MAXIGP1AWID(pps$MAXIGP1AWID),
        .MAXIGP1AWLEN(pps$MAXIGP1AWLEN),
        .MAXIGP1AWLOCK(pps$MAXIGP1AWLOCK),
        .MAXIGP1AWPROT(pps$MAXIGP1AWPROT),
        .MAXIGP1AWQOS(pps$MAXIGP1AWQOS),
        .MAXIGP1AWREADY(pps$MAXIGP1AWREADY),
        .MAXIGP1AWSIZE(pps$MAXIGP1AWSIZE),
        .MAXIGP1AWVALID(pps$MAXIGP1AWVALID),
        .MAXIGP1BID(pps$MAXIGP1BID),
        .MAXIGP1BREADY(pps$MAXIGP1BREADY),
        .MAXIGP1BRESP(pps$MAXIGP1BRESP),
        .MAXIGP1BVALID(pps$MAXIGP1BVALID),
        .MAXIGP1RDATA(pps$MAXIGP1RDATA),
        .MAXIGP1RID(pps$MAXIGP1RID),
        .MAXIGP1RLAST(pps$MAXIGP1RLAST),
        .MAXIGP1RREADY(pps$MAXIGP1RREADY),
        .MAXIGP1RRESP(pps$MAXIGP1RRESP),
        .MAXIGP1RVALID(pps$MAXIGP1RVALID),
        .MAXIGP1WDATA(pps$MAXIGP1WDATA),
        .MAXIGP1WID(pps$MAXIGP1WID),
        .MAXIGP1WLAST(pps$MAXIGP1WLAST),
        .MAXIGP1WREADY(pps$MAXIGP1WREADY),
        .MAXIGP1WSTRB(pps$MAXIGP1WSTRB),
        .MAXIGP1WVALID(pps$MAXIGP1WVALID),
        .MIO(MIO),
        .PSCLK(PSCLK),
        .PSPORB(PSPORB),
        .PSSRSTB(PSSRSTB),
        .SAXIACPACLK(CLK),
        .SAXIACPARADDR(pps$SAXIACPARADDR),
        .SAXIACPARBURST(pps$SAXIACPARBURST),
        .SAXIACPARCACHE(pps$SAXIACPARCACHE),
        .SAXIACPARESETN(pps$SAXIACPARESETN),
        .SAXIACPARID(pps$SAXIACPARID),
        .SAXIACPARLEN(pps$SAXIACPARLEN),
        .SAXIACPARLOCK(pps$SAXIACPARLOCK),
        .SAXIACPARPROT(pps$SAXIACPARPROT),
        .SAXIACPARQOS(pps$SAXIACPARQOS),
        .SAXIACPARREADY(pps$SAXIACPARREADY),
        .SAXIACPARSIZE(pps$SAXIACPARSIZE),
        .SAXIACPARUSER(pps$SAXIACPARUSER),
        .SAXIACPARVALID(pps$SAXIACPARVALID),
        .SAXIACPAWADDR(pps$SAXIACPAWADDR),
        .SAXIACPAWBURST(pps$SAXIACPAWBURST),
        .SAXIACPAWCACHE(pps$SAXIACPAWCACHE),
        .SAXIACPAWID(pps$SAXIACPAWID),
        .SAXIACPAWLEN(pps$SAXIACPAWLEN),
        .SAXIACPAWLOCK(pps$SAXIACPAWLOCK),
        .SAXIACPAWPROT(pps$SAXIACPAWPROT),
        .SAXIACPAWQOS(pps$SAXIACPAWQOS),
        .SAXIACPAWREADY(pps$SAXIACPAWREADY),
        .SAXIACPAWSIZE(pps$SAXIACPAWSIZE),
        .SAXIACPAWUSER(pps$SAXIACPAWUSER),
        .SAXIACPAWVALID(pps$SAXIACPAWVALID),
        .SAXIACPBID(pps$SAXIACPBID),
        .SAXIACPBREADY(pps$SAXIACPBREADY),
        .SAXIACPBRESP(pps$SAXIACPBRESP),
        .SAXIACPBVALID(pps$SAXIACPBVALID),
        .SAXIACPRDATA(pps$SAXIACPRDATA),
        .SAXIACPRID(pps$SAXIACPRID),
        .SAXIACPRLAST(pps$SAXIACPRLAST),
        .SAXIACPRREADY(pps$SAXIACPRREADY),
        .SAXIACPRRESP(pps$SAXIACPRRESP),
        .SAXIACPRVALID(pps$SAXIACPRVALID),
        .SAXIACPWDATA(pps$SAXIACPWDATA),
        .SAXIACPWID(pps$SAXIACPWID),
        .SAXIACPWLAST(pps$SAXIACPWLAST),
        .SAXIACPWREADY(pps$SAXIACPWREADY),
        .SAXIACPWSTRB(pps$SAXIACPWSTRB),
        .SAXIACPWVALID(pps$SAXIACPWVALID),
        .SAXIGP0ACLK(CLK),
        .SAXIGP0ARADDR(pps$SAXIGP0ARADDR),
        .SAXIGP0ARBURST(pps$SAXIGP0ARBURST),
        .SAXIGP0ARCACHE(pps$SAXIGP0ARCACHE),
        .SAXIGP0ARESETN(pps$SAXIGP0ARESETN),
        .SAXIGP0ARID(pps$SAXIGP0ARID),
        .SAXIGP0ARLEN(pps$SAXIGP0ARLEN),
        .SAXIGP0ARLOCK(pps$SAXIGP0ARLOCK),
        .SAXIGP0ARPROT(pps$SAXIGP0ARPROT),
        .SAXIGP0ARQOS(pps$SAXIGP0ARQOS),
        .SAXIGP0ARREADY(pps$SAXIGP0ARREADY),
        .SAXIGP0ARSIZE(pps$SAXIGP0ARSIZE),
        .SAXIGP0ARVALID(pps$SAXIGP0ARVALID),
        .SAXIGP0AWADDR(pps$SAXIGP0AWADDR),
        .SAXIGP0AWBURST(pps$SAXIGP0AWBURST),
        .SAXIGP0AWCACHE(pps$SAXIGP0AWCACHE),
        .SAXIGP0AWID(pps$SAXIGP0AWID),
        .SAXIGP0AWLEN(pps$SAXIGP0AWLEN),
        .SAXIGP0AWLOCK(pps$SAXIGP0AWLOCK),
        .SAXIGP0AWPROT(pps$SAXIGP0AWPROT),
        .SAXIGP0AWQOS(pps$SAXIGP0AWQOS),
        .SAXIGP0AWREADY(pps$SAXIGP0AWREADY),
        .SAXIGP0AWSIZE(pps$SAXIGP0AWSIZE),
        .SAXIGP0AWVALID(pps$SAXIGP0AWVALID),
        .SAXIGP0BID(pps$SAXIGP0BID),
        .SAXIGP0BREADY(pps$SAXIGP0BREADY),
        .SAXIGP0BRESP(pps$SAXIGP0BRESP),
        .SAXIGP0BVALID(pps$SAXIGP0BVALID),
        .SAXIGP0RDATA(pps$SAXIGP0RDATA),
        .SAXIGP0RID(pps$SAXIGP0RID),
        .SAXIGP0RLAST(pps$SAXIGP0RLAST),
        .SAXIGP0RREADY(pps$SAXIGP0RREADY),
        .SAXIGP0RRESP(pps$SAXIGP0RRESP),
        .SAXIGP0RVALID(pps$SAXIGP0RVALID),
        .SAXIGP0WDATA(pps$SAXIGP0WDATA),
        .SAXIGP0WID(pps$SAXIGP0WID),
        .SAXIGP0WLAST(pps$SAXIGP0WLAST),
        .SAXIGP0WREADY(pps$SAXIGP0WREADY),
        .SAXIGP0WSTRB(pps$SAXIGP0WSTRB),
        .SAXIGP0WVALID(pps$SAXIGP0WVALID),
        .SAXIGP1ACLK(CLK),
        .SAXIGP1ARADDR(pps$SAXIGP1ARADDR),
        .SAXIGP1ARBURST(pps$SAXIGP1ARBURST),
        .SAXIGP1ARCACHE(pps$SAXIGP1ARCACHE),
        .SAXIGP1ARESETN(pps$SAXIGP1ARESETN),
        .SAXIGP1ARID(pps$SAXIGP1ARID),
        .SAXIGP1ARLEN(pps$SAXIGP1ARLEN),
        .SAXIGP1ARLOCK(pps$SAXIGP1ARLOCK),
        .SAXIGP1ARPROT(pps$SAXIGP1ARPROT),
        .SAXIGP1ARQOS(pps$SAXIGP1ARQOS),
        .SAXIGP1ARREADY(pps$SAXIGP1ARREADY),
        .SAXIGP1ARSIZE(pps$SAXIGP1ARSIZE),
        .SAXIGP1ARVALID(pps$SAXIGP1ARVALID),
        .SAXIGP1AWADDR(pps$SAXIGP1AWADDR),
        .SAXIGP1AWBURST(pps$SAXIGP1AWBURST),
        .SAXIGP1AWCACHE(pps$SAXIGP1AWCACHE),
        .SAXIGP1AWID(pps$SAXIGP1AWID),
        .SAXIGP1AWLEN(pps$SAXIGP1AWLEN),
        .SAXIGP1AWLOCK(pps$SAXIGP1AWLOCK),
        .SAXIGP1AWPROT(pps$SAXIGP1AWPROT),
        .SAXIGP1AWQOS(pps$SAXIGP1AWQOS),
        .SAXIGP1AWREADY(pps$SAXIGP1AWREADY),
        .SAXIGP1AWSIZE(pps$SAXIGP1AWSIZE),
        .SAXIGP1AWVALID(pps$SAXIGP1AWVALID),
        .SAXIGP1BID(pps$SAXIGP1BID),
        .SAXIGP1BREADY(pps$SAXIGP1BREADY),
        .SAXIGP1BRESP(pps$SAXIGP1BRESP),
        .SAXIGP1BVALID(pps$SAXIGP1BVALID),
        .SAXIGP1RDATA(pps$SAXIGP1RDATA),
        .SAXIGP1RID(pps$SAXIGP1RID),
        .SAXIGP1RLAST(pps$SAXIGP1RLAST),
        .SAXIGP1RREADY(pps$SAXIGP1RREADY),
        .SAXIGP1RRESP(pps$SAXIGP1RRESP),
        .SAXIGP1RVALID(pps$SAXIGP1RVALID),
        .SAXIGP1WDATA(pps$SAXIGP1WDATA),
        .SAXIGP1WID(pps$SAXIGP1WID),
        .SAXIGP1WLAST(pps$SAXIGP1WLAST),
        .SAXIGP1WREADY(pps$SAXIGP1WREADY),
        .SAXIGP1WSTRB(pps$SAXIGP1WSTRB),
        .SAXIGP1WVALID(pps$SAXIGP1WVALID),
        .SAXIHP0ACLK(CLK),
        .SAXIHP0ARADDR(pps$SAXIHP0ARADDR),
        .SAXIHP0ARBURST(pps$SAXIHP0ARBURST),
        .SAXIHP0ARCACHE(pps$SAXIHP0ARCACHE),
        .SAXIHP0ARESETN(pps$SAXIHP0ARESETN),
        .SAXIHP0ARID(pps$SAXIHP0ARID),
        .SAXIHP0ARLEN(pps$SAXIHP0ARLEN),
        .SAXIHP0ARLOCK(pps$SAXIHP0ARLOCK),
        .SAXIHP0ARPROT(pps$SAXIHP0ARPROT),
        .SAXIHP0ARQOS(pps$SAXIHP0ARQOS),
        .SAXIHP0ARREADY(pps$SAXIHP0ARREADY),
        .SAXIHP0ARSIZE(pps$SAXIHP0ARSIZE),
        .SAXIHP0ARVALID(pps$SAXIHP0ARVALID),
        .SAXIHP0AWADDR(pps$SAXIHP0AWADDR),
        .SAXIHP0AWBURST(pps$SAXIHP0AWBURST),
        .SAXIHP0AWCACHE(pps$SAXIHP0AWCACHE),
        .SAXIHP0AWID(pps$SAXIHP0AWID),
        .SAXIHP0AWLEN(pps$SAXIHP0AWLEN),
        .SAXIHP0AWLOCK(pps$SAXIHP0AWLOCK),
        .SAXIHP0AWPROT(pps$SAXIHP0AWPROT),
        .SAXIHP0AWQOS(pps$SAXIHP0AWQOS),
        .SAXIHP0AWREADY(pps$SAXIHP0AWREADY),
        .SAXIHP0AWSIZE(pps$SAXIHP0AWSIZE),
        .SAXIHP0AWVALID(pps$SAXIHP0AWVALID),
        .SAXIHP0BID(pps$SAXIHP0BID),
        .SAXIHP0BREADY(pps$SAXIHP0BREADY),
        .SAXIHP0BRESP(pps$SAXIHP0BRESP),
        .SAXIHP0BVALID(pps$SAXIHP0BVALID),
        .SAXIHP0RACOUNT(pps$SAXIHP0RACOUNT),
        .SAXIHP0RCOUNT(pps$SAXIHP0RCOUNT),
        .SAXIHP0RDATA(pps$SAXIHP0RDATA),
        .SAXIHP0RDISSUECAP1EN(pps$SAXIHP0RDISSUECAP1EN),
        .SAXIHP0RID(pps$SAXIHP0RID),
        .SAXIHP0RLAST(pps$SAXIHP0RLAST),
        .SAXIHP0RREADY(pps$SAXIHP0RREADY),
        .SAXIHP0RRESP(pps$SAXIHP0RRESP),
        .SAXIHP0RVALID(pps$SAXIHP0RVALID),
        .SAXIHP0WACOUNT(pps$SAXIHP0WACOUNT),
        .SAXIHP0WCOUNT(pps$SAXIHP0WCOUNT),
        .SAXIHP0WDATA(pps$SAXIHP0WDATA),
        .SAXIHP0WID(pps$SAXIHP0WID),
        .SAXIHP0WLAST(pps$SAXIHP0WLAST),
        .SAXIHP0WREADY(pps$SAXIHP0WREADY),
        .SAXIHP0WRISSUECAP1EN(pps$SAXIHP0WRISSUECAP1EN),
        .SAXIHP0WSTRB(pps$SAXIHP0WSTRB),
        .SAXIHP0WVALID(pps$SAXIHP0WVALID),
        .SAXIHP1ACLK(CLK),
        .SAXIHP1ARADDR(pps$SAXIHP1ARADDR),
        .SAXIHP1ARBURST(pps$SAXIHP1ARBURST),
        .SAXIHP1ARCACHE(pps$SAXIHP1ARCACHE),
        .SAXIHP1ARESETN(pps$SAXIHP1ARESETN),
        .SAXIHP1ARID(pps$SAXIHP1ARID),
        .SAXIHP1ARLEN(pps$SAXIHP1ARLEN),
        .SAXIHP1ARLOCK(pps$SAXIHP1ARLOCK),
        .SAXIHP1ARPROT(pps$SAXIHP1ARPROT),
        .SAXIHP1ARQOS(pps$SAXIHP1ARQOS),
        .SAXIHP1ARREADY(pps$SAXIHP1ARREADY),
        .SAXIHP1ARSIZE(pps$SAXIHP1ARSIZE),
        .SAXIHP1ARVALID(pps$SAXIHP1ARVALID),
        .SAXIHP1AWADDR(pps$SAXIHP1AWADDR),
        .SAXIHP1AWBURST(pps$SAXIHP1AWBURST),
        .SAXIHP1AWCACHE(pps$SAXIHP1AWCACHE),
        .SAXIHP1AWID(pps$SAXIHP1AWID),
        .SAXIHP1AWLEN(pps$SAXIHP1AWLEN),
        .SAXIHP1AWLOCK(pps$SAXIHP1AWLOCK),
        .SAXIHP1AWPROT(pps$SAXIHP1AWPROT),
        .SAXIHP1AWQOS(pps$SAXIHP1AWQOS),
        .SAXIHP1AWREADY(pps$SAXIHP1AWREADY),
        .SAXIHP1AWSIZE(pps$SAXIHP1AWSIZE),
        .SAXIHP1AWVALID(pps$SAXIHP1AWVALID),
        .SAXIHP1BID(pps$SAXIHP1BID),
        .SAXIHP1BREADY(pps$SAXIHP1BREADY),
        .SAXIHP1BRESP(pps$SAXIHP1BRESP),
        .SAXIHP1BVALID(pps$SAXIHP1BVALID),
        .SAXIHP1RACOUNT(pps$SAXIHP1RACOUNT),
        .SAXIHP1RCOUNT(pps$SAXIHP1RCOUNT),
        .SAXIHP1RDATA(pps$SAXIHP1RDATA),
        .SAXIHP1RDISSUECAP1EN(pps$SAXIHP1RDISSUECAP1EN),
        .SAXIHP1RID(pps$SAXIHP1RID),
        .SAXIHP1RLAST(pps$SAXIHP1RLAST),
        .SAXIHP1RREADY(pps$SAXIHP1RREADY),
        .SAXIHP1RRESP(pps$SAXIHP1RRESP),
        .SAXIHP1RVALID(pps$SAXIHP1RVALID),
        .SAXIHP1WACOUNT(pps$SAXIHP1WACOUNT),
        .SAXIHP1WCOUNT(pps$SAXIHP1WCOUNT),
        .SAXIHP1WDATA(pps$SAXIHP1WDATA),
        .SAXIHP1WID(pps$SAXIHP1WID),
        .SAXIHP1WLAST(pps$SAXIHP1WLAST),
        .SAXIHP1WREADY(pps$SAXIHP1WREADY),
        .SAXIHP1WRISSUECAP1EN(pps$SAXIHP1WRISSUECAP1EN),
        .SAXIHP1WSTRB(pps$SAXIHP1WSTRB),
        .SAXIHP1WVALID(pps$SAXIHP1WVALID),
        .SAXIHP2ACLK(CLK),
        .SAXIHP2ARADDR(pps$SAXIHP2ARADDR),
        .SAXIHP2ARBURST(pps$SAXIHP2ARBURST),
        .SAXIHP2ARCACHE(pps$SAXIHP2ARCACHE),
        .SAXIHP2ARESETN(pps$SAXIHP2ARESETN),
        .SAXIHP2ARID(pps$SAXIHP2ARID),
        .SAXIHP2ARLEN(pps$SAXIHP2ARLEN),
        .SAXIHP2ARLOCK(pps$SAXIHP2ARLOCK),
        .SAXIHP2ARPROT(pps$SAXIHP2ARPROT),
        .SAXIHP2ARQOS(pps$SAXIHP2ARQOS),
        .SAXIHP2ARREADY(pps$SAXIHP2ARREADY),
        .SAXIHP2ARSIZE(pps$SAXIHP2ARSIZE),
        .SAXIHP2ARVALID(pps$SAXIHP2ARVALID),
        .SAXIHP2AWADDR(pps$SAXIHP2AWADDR),
        .SAXIHP2AWBURST(pps$SAXIHP2AWBURST),
        .SAXIHP2AWCACHE(pps$SAXIHP2AWCACHE),
        .SAXIHP2AWID(pps$SAXIHP2AWID),
        .SAXIHP2AWLEN(pps$SAXIHP2AWLEN),
        .SAXIHP2AWLOCK(pps$SAXIHP2AWLOCK),
        .SAXIHP2AWPROT(pps$SAXIHP2AWPROT),
        .SAXIHP2AWQOS(pps$SAXIHP2AWQOS),
        .SAXIHP2AWREADY(pps$SAXIHP2AWREADY),
        .SAXIHP2AWSIZE(pps$SAXIHP2AWSIZE),
        .SAXIHP2AWVALID(pps$SAXIHP2AWVALID),
        .SAXIHP2BID(pps$SAXIHP2BID),
        .SAXIHP2BREADY(pps$SAXIHP2BREADY),
        .SAXIHP2BRESP(pps$SAXIHP2BRESP),
        .SAXIHP2BVALID(pps$SAXIHP2BVALID),
        .SAXIHP2RACOUNT(pps$SAXIHP2RACOUNT),
        .SAXIHP2RCOUNT(pps$SAXIHP2RCOUNT),
        .SAXIHP2RDATA(pps$SAXIHP2RDATA),
        .SAXIHP2RDISSUECAP1EN(pps$SAXIHP2RDISSUECAP1EN),
        .SAXIHP2RID(pps$SAXIHP2RID),
        .SAXIHP2RLAST(pps$SAXIHP2RLAST),
        .SAXIHP2RREADY(pps$SAXIHP2RREADY),
        .SAXIHP2RRESP(pps$SAXIHP2RRESP),
        .SAXIHP2RVALID(pps$SAXIHP2RVALID),
        .SAXIHP2WACOUNT(pps$SAXIHP2WACOUNT),
        .SAXIHP2WCOUNT(pps$SAXIHP2WCOUNT),
        .SAXIHP2WDATA(pps$SAXIHP2WDATA),
        .SAXIHP2WID(pps$SAXIHP2WID),
        .SAXIHP2WLAST(pps$SAXIHP2WLAST),
        .SAXIHP2WREADY(pps$SAXIHP2WREADY),
        .SAXIHP2WRISSUECAP1EN(pps$SAXIHP2WRISSUECAP1EN),
        .SAXIHP2WSTRB(pps$SAXIHP2WSTRB),
        .SAXIHP2WVALID(pps$SAXIHP2WVALID),
        .SAXIHP3ACLK(CLK),
        .SAXIHP3ARADDR(pps$SAXIHP3ARADDR),
        .SAXIHP3ARBURST(pps$SAXIHP3ARBURST),
        .SAXIHP3ARCACHE(pps$SAXIHP3ARCACHE),
        .SAXIHP3ARESETN(pps$SAXIHP3ARESETN),
        .SAXIHP3ARID(pps$SAXIHP3ARID),
        .SAXIHP3ARLEN(pps$SAXIHP3ARLEN),
        .SAXIHP3ARLOCK(pps$SAXIHP3ARLOCK),
        .SAXIHP3ARPROT(pps$SAXIHP3ARPROT),
        .SAXIHP3ARQOS(pps$SAXIHP3ARQOS),
        .SAXIHP3ARREADY(pps$SAXIHP3ARREADY),
        .SAXIHP3ARSIZE(pps$SAXIHP3ARSIZE),
        .SAXIHP3ARVALID(pps$SAXIHP3ARVALID),
        .SAXIHP3AWADDR(pps$SAXIHP3AWADDR),
        .SAXIHP3AWBURST(pps$SAXIHP3AWBURST),
        .SAXIHP3AWCACHE(pps$SAXIHP3AWCACHE),
        .SAXIHP3AWID(pps$SAXIHP3AWID),
        .SAXIHP3AWLEN(pps$SAXIHP3AWLEN),
        .SAXIHP3AWLOCK(pps$SAXIHP3AWLOCK),
        .SAXIHP3AWPROT(pps$SAXIHP3AWPROT),
        .SAXIHP3AWQOS(pps$SAXIHP3AWQOS),
        .SAXIHP3AWREADY(pps$SAXIHP3AWREADY),
        .SAXIHP3AWSIZE(pps$SAXIHP3AWSIZE),
        .SAXIHP3AWVALID(pps$SAXIHP3AWVALID),
        .SAXIHP3BID(pps$SAXIHP3BID),
        .SAXIHP3BREADY(pps$SAXIHP3BREADY),
        .SAXIHP3BRESP(pps$SAXIHP3BRESP),
        .SAXIHP3BVALID(pps$SAXIHP3BVALID),
        .SAXIHP3RACOUNT(pps$SAXIHP3RACOUNT),
        .SAXIHP3RCOUNT(pps$SAXIHP3RCOUNT),
        .SAXIHP3RDATA(pps$SAXIHP3RDATA),
        .SAXIHP3RDISSUECAP1EN(pps$SAXIHP3RDISSUECAP1EN),
        .SAXIHP3RID(pps$SAXIHP3RID),
        .SAXIHP3RLAST(pps$SAXIHP3RLAST),
        .SAXIHP3RREADY(pps$SAXIHP3RREADY),
        .SAXIHP3RRESP(pps$SAXIHP3RRESP),
        .SAXIHP3RVALID(pps$SAXIHP3RVALID),
        .SAXIHP3WACOUNT(pps$SAXIHP3WACOUNT),
        .SAXIHP3WCOUNT(pps$SAXIHP3WCOUNT),
        .SAXIHP3WDATA(pps$SAXIHP3WDATA),
        .SAXIHP3WID(pps$SAXIHP3WID),
        .SAXIHP3WLAST(pps$SAXIHP3WLAST),
        .SAXIHP3WREADY(pps$SAXIHP3WREADY),
        .SAXIHP3WRISSUECAP1EN(pps$SAXIHP3WRISSUECAP1EN),
        .SAXIHP3WSTRB(pps$SAXIHP3WSTRB),
        .SAXIHP3WVALID(pps$SAXIHP3WVALID));
    BUFG ps7_fclk_0_c (
        .I(FCLKCLK),
        .O(CLK));
    BUFG ps7_freset_0_r (
        .I(pps$FCLKRESETN),
        .O(nRST));
    assign pps$DMA0ACLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA0DAREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA0DRLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA0DRTYPE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA0DRVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA1ACLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA1DAREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA1DRLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA1DRTYPE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA1DRVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA2ACLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA2DAREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA2DRLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA2DRTYPE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA2DRVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA3ACLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA3DAREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA3DRLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA3DRTYPE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$DMA3DRVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOCAN0PHYRX = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOCAN1PHYRX = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0EXTINTIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIICOL = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIICRS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIIRXCLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIIRXD = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIIRXDV = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIIRXER = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0GMIITXCLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET0MDIOI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1EXTINTIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIICOL = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIICRS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIIRXCLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIIRXD = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIIRXDV = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIIRXER = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1GMIITXCLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOENET1MDIOI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOGPIOI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOI2C0SCLI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOI2C0SDAI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOI2C1SCLI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOI2C1SDAI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOPJTAGTCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOPJTAGTDI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOPJTAGTMS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO0CDN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO0CLKFB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO0CMDI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO0DATAI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO0WP = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO1CDN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO1CLKFB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO1CMDI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO1DATAI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSDIO1WP = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI0MI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI0SCLKI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI0SI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI0SSIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI1MI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI1SCLKI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI1SI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSPI1SSIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOSRAMINTIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOTRACECLK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOTTC0CLKI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOTTC1CLKI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART0CTSN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART0DCDN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART0DSRN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART0RIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART0RX = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART1CTSN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART1DCDN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART1DSRN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART1RIN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUART1RX = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUSB0VBUSPWRFAULT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOUSB1VBUSPWRFAULT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EMIOWDTCLKI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$EVENTEVENTI = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FCLKCLKTRIGN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMDTRACEINATID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMDTRACEINCLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMDTRACEINDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMDTRACEINVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMTF2PDEBUG = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMTF2PTRIG = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$FTMTP2FTRIGACK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1ARREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1AWREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1BID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1BRESP = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1BVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1RDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1RID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1RLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1RRESP = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1RVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$MAXIGP1WREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARUSER = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWUSER = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPAWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPBREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPRREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPWDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPWLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPWSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIACPWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP0WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIGP1WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0RDISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WRISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP0WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1RDISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WRISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP1WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2RDISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WRISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP2WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3ARVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWADDR = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWBURST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWCACHE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWLEN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWLOCK = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWPROT = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWQOS = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWSIZE = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3AWVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3BREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3RDISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3RREADY = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WDATA = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WLAST = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WRISSUECAP1EN = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WSTRB = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
    assign pps$SAXIHP3WVALID = 0; //MISSING_ASSIGNMENT_FOR_OUTPUT_VALUE
endmodule 

