`ifndef __mimo_GENERATED__VH__
`define __mimo_GENERATED__VH__

//METASTART; MIMOBase
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; !( c >= widthOut );
//METAGUARD; out$deq; c >= widthOut;
//METAGUARD; out$first; c >= widthOut;
`endif
