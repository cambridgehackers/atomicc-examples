`include "atomicclib.vh"

//METASTART; SyncFF
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$init
