`ifndef __printfStub_GENERATED__VH__
`define __printfStub_GENERATED__VH__
`include "atomicclib.vh"

//METASTART; Printf
//METAGUARD; enq; 1'd1;
`endif
