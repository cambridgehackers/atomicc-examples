`ifndef __iobufVec_GENERATED__VH__
`define __iobufVec_GENERATED__VH__

//METASTART; IobufVec
//METAINTERNAL; iobufs0; IOBUF;
//METAGUARD; RULE$iobufs; 1'd1;
//METARULES; RULE$iobufs
`endif
