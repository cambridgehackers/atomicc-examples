`ifndef __vsimTop_GENERATED__VH__
`define __vsimTop_GENERATED__VH__

//METASTART; VsimTop
//METAINTERNAL; user; UserTop;
//METAINTERNAL; sink_0; VsimReceive(width=32);
//METAINTERNAL; source_0; VsimSend(width=32);
//METACONNECT; sink_0$$enq__ENA; user$write$enq__ENA
//METACONNECT; sink_0$$enq__RDY; user$write$enq__RDY
//METACONNECT; user$read$enq__ENA; source_0$enq__ENA
//METACONNECT; user$read$enq__RDY; source_0$enq__RDY
`endif
