`ifndef __funnel_GENERATED__VH__
`define __funnel_GENERATED__VH__

//METASTART; FunnelHalfBase
//METAEXTERNAL; output; FunnelHalfBase$output;
//METAGUARD; input$enq; ( ( ( ( __inst$Genvar1 + 1 ) / 2 ) == ( __inst$Genvar1 / 2 ) ) && ( output[ __inst$Genvar1 / 2 ] . enq__RDY ) ) || ( ( !( ( ( __inst$Genvar1 + 1 ) / 2 ) == ( __inst$Genvar1 / 2 ) ) ) && ( output[ __inst$Genvar1 / 2 ] . enq__RDY ) && ( enq__ENA == 0 ) );
`endif
