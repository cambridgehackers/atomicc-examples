`ifndef __printfStub_GENERATED__VH__
`define __printfStub_GENERATED__VH__

//METASTART; Printf
//METAGUARD; enq; 1;
`endif
