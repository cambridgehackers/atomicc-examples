`ifndef __gearNto1_GENERATED__VH__
`define __gearNto1_GENERATED__VH__

//METASTART; GearNto1Base
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; c == 0;
//METAGUARD; out$deq; !( c == 0 );
//METAGUARD; out$first; !( c == 0 );
`endif
