`include "ivector.generated.vh"

module l_module_OC_Fifo1 (
    input CLK,
    input nRST,
    input out$deq__ENA,
    output out$deq__RDY,
    input in$enq__ENA,
    input [31:0]in$enq_v,
    output in$enq__RDY,
    output [31:0]out$first,
    output out$first__RDY);
    wire out$deq__RDY_internal;
    wire out$deq__ENA_internal = out$deq__ENA && out$deq__RDY_internal;
    wire in$enq__RDY_internal;
    wire in$enq__ENA_internal = in$enq__ENA && in$enq__RDY_internal;
    reg[31:0] element;
    reg full;
    assign in$enq__RDY = in$enq__RDY_internal;
    assign in$enq__RDY_internal = full ^ 1;
    assign out$deq__RDY = out$deq__RDY_internal;
    assign out$deq__RDY_internal = full;
    assign out$first = element;
    assign out$first__RDY_internal = full;

    always @( posedge CLK) begin
      if (!nRST) begin
        element <= 0;
        full <= 0;
      end // nRST
      else begin
        if (out$deq__ENA_internal) begin
            full <= 0;
        end; // End of out$deq__ENA
        if (in$enq__ENA_internal) begin
            element <= in$enq_v;
            full <= 1;
        end; // End of in$enq__ENA
      end
    end // always @ (posedge CLK)
endmodule 

module l_module_OC_Fifo1_OC_3 (
    input CLK,
    input nRST,
    input out$deq__ENA,
    output out$deq__RDY,
    input in$enq__ENA,
    input [95:0]in$enq_v,
    output in$enq__RDY,
    output [95:0]out$first,
    output out$first__RDY);
    wire out$deq__RDY_internal;
    wire out$deq__ENA_internal = out$deq__ENA && out$deq__RDY_internal;
    wire in$enq__RDY_internal;
    wire in$enq__ENA_internal = in$enq__ENA && in$enq__RDY_internal;
    reg[95:0] element;
    reg full;
    assign in$enq__RDY = in$enq__RDY_internal;
    assign in$enq__RDY_internal = full ^ 1;
    assign out$deq__RDY = out$deq__RDY_internal;
    assign out$deq__RDY_internal = full;
    assign out$first = element;
    assign out$first__RDY_internal = full;

    always @( posedge CLK) begin
      if (!nRST) begin
        element <= 0;
        full <= 0;
      end // nRST
      else begin
        if (out$deq__ENA_internal) begin
            full <= 0;
        end; // End of out$deq__ENA
        if (in$enq__ENA_internal) begin
            element <= in$enq_v;
            full <= 1;
        end; // End of in$enq__ENA
      end
    end // always @ (posedge CLK)
endmodule 

module l_module_OC_FifoPong (
    input CLK,
    input nRST,
    input out$deq__ENA,
    output out$deq__RDY,
    input in$enq__ENA,
    input [95:0]in$enq_v,
    output in$enq__RDY,
    output [95:0]out$first,
    output out$first__RDY);
    wire out$deq__RDY_internal;
    wire out$deq__ENA_internal = out$deq__ENA && out$deq__RDY_internal;
    wire in$enq__RDY_internal;
    wire in$enq__ENA_internal = in$enq__ENA && in$enq__RDY_internal;
    wire element1$out$deq__RDY;
    wire element1$in$enq__RDY;
    wire [95:0]element1$out$first;
    wire element1$out$first__RDY;
    l_module_OC_Fifo1_OC_3 element1 (
        CLK,
        nRST,
        out$deq__ENA_internal & pong ^ 1,
        element1$out$deq__RDY,
        in$enq__ENA_internal & pong ^ 1,
        element2$in$enq_v,
        element1$in$enq__RDY,
        element1$out$first,
        element1$out$first__RDY);
    wire element2$out$deq__RDY;
    wire [95:0]element2$in$enq_v;
    wire element2$in$enq__RDY;
    wire [95:0]element2$out$first;
    wire element2$out$first__RDY;
    l_module_OC_Fifo1_OC_3 element2 (
        CLK,
        nRST,
        out$deq__ENA_internal & pong,
        element2$out$deq__RDY,
        in$enq__ENA_internal & pong,
        element2$in$enq_v,
        element2$in$enq__RDY,
        element2$out$first,
        element2$out$first__RDY);
    reg pong;
    assign in$enq__RDY = in$enq__RDY_internal;
    assign in$enq__RDY_internal = (element2$in$enq__RDY | (pong ^ 1)) & (element1$in$enq__RDY | pong);
    assign out$deq__RDY = out$deq__RDY_internal;
    assign out$deq__RDY_internal = (element2$out$deq__RDY | (pong ^ 1)) & (element1$out$deq__RDY | pong);
    assign out$first = retval;
    assign out$first__RDY_internal = (element2$out$first__RDY | (pong ^ 1)) & (element1$out$first__RDY | pong);
    assign retval$a = element1$out$first.a;
    assign retval$b = element1$out$first.b;
    assign retval$c = element1$out$first.c;

    always @( posedge CLK) begin
      if (!nRST) begin
        pong <= 0;
      end // nRST
      else begin
        if (out$deq__ENA_internal) begin
            pong <= pong ^ 1;
        end; // End of out$deq__ENA
      end
    end // always @ (posedge CLK)
endmodule 

module l_module_OC_IVector (
    input CLK,
    input nRST,
    input in$say__ENA,
    input [31:0]in$say_meth,
    input [31:0]in$say_v,
    output in$say__RDY,
    output ind$heard__ENA,
    output [31:0]ind$heard_heard_meth,
    output [31:0]ind$heard_heard_v,
    input ind$heard__RDY);
    wire in$say__RDY_internal;
    wire in$say__ENA_internal = in$say__ENA && in$say__RDY_internal;
    wire fifo0$out$deq__RDY;
    wire fifo0$in$enq__ENA;
    wire [95:0]fifo0$in$enq_v;
    wire fifo0$in$enq__RDY;
    wire [95:0]fifo0$out$first;
    wire fifo0$out$first__RDY;
    l_module_OC_FifoPong fifo0 (
        CLK,
        nRST,
        respond0__ENA_internal,
        fifo0$out$deq__RDY,
        fifo0$in$enq__ENA,
        fifo0$in$enq_v,
        fifo0$in$enq__RDY,
        fifo0$out$first,
        fifo0$out$first__RDY);
    wire fifo1$out$deq__RDY;
    wire fifo1$in$enq__ENA;
    wire [95:0]fifo1$in$enq_v;
    wire fifo1$in$enq__RDY;
    wire [95:0]fifo1$out$first;
    wire fifo1$out$first__RDY;
    l_module_OC_FifoPong fifo1 (
        CLK,
        nRST,
        respond1__ENA_internal,
        fifo1$out$deq__RDY,
        fifo1$in$enq__ENA,
        fifo1$in$enq_v,
        fifo1$in$enq__RDY,
        fifo1$out$first,
        fifo1$out$first__RDY);
    wire fifo2$out$deq__RDY;
    wire fifo2$in$enq__ENA;
    wire [95:0]fifo2$in$enq_v;
    wire fifo2$in$enq__RDY;
    wire [95:0]fifo2$out$first;
    wire fifo2$out$first__RDY;
    l_module_OC_FifoPong fifo2 (
        CLK,
        nRST,
        respond2__ENA_internal,
        fifo2$out$deq__RDY,
        fifo2$in$enq__ENA,
        fifo2$in$enq_v,
        fifo2$in$enq__RDY,
        fifo2$out$first,
        fifo2$out$first__RDY);
    wire fifo3$out$deq__RDY;
    wire fifo3$in$enq__ENA;
    wire [95:0]fifo3$in$enq_v;
    wire fifo3$in$enq__RDY;
    wire [95:0]fifo3$out$first;
    wire fifo3$out$first__RDY;
    l_module_OC_FifoPong fifo3 (
        CLK,
        nRST,
        respond3__ENA_internal,
        fifo3$out$deq__RDY,
        fifo3$in$enq__ENA,
        fifo3$in$enq_v,
        fifo3$in$enq__RDY,
        fifo3$out$first,
        fifo3$out$first__RDY);
    wire fifo4$out$deq__RDY;
    wire fifo4$in$enq__ENA;
    wire [95:0]fifo4$in$enq_v;
    wire fifo4$in$enq__RDY;
    wire [95:0]fifo4$out$first;
    wire fifo4$out$first__RDY;
    l_module_OC_FifoPong fifo4 (
        CLK,
        nRST,
        respond4__ENA_internal,
        fifo4$out$deq__RDY,
        fifo4$in$enq__ENA,
        fifo4$in$enq_v,
        fifo4$in$enq__RDY,
        fifo4$out$first,
        fifo4$out$first__RDY);
    wire fifo5$out$deq__RDY;
    wire fifo5$in$enq__ENA;
    wire [95:0]fifo5$in$enq_v;
    wire fifo5$in$enq__RDY;
    wire [95:0]fifo5$out$first;
    wire fifo5$out$first__RDY;
    l_module_OC_FifoPong fifo5 (
        CLK,
        nRST,
        respond5__ENA_internal,
        fifo5$out$deq__RDY,
        fifo5$in$enq__ENA,
        fifo5$in$enq_v,
        fifo5$in$enq__RDY,
        fifo5$out$first,
        fifo5$out$first__RDY);
    wire fifo6$out$deq__RDY;
    wire fifo6$in$enq__ENA;
    wire [95:0]fifo6$in$enq_v;
    wire fifo6$in$enq__RDY;
    wire [95:0]fifo6$out$first;
    wire fifo6$out$first__RDY;
    l_module_OC_FifoPong fifo6 (
        CLK,
        nRST,
        respond6__ENA_internal,
        fifo6$out$deq__RDY,
        fifo6$in$enq__ENA,
        fifo6$in$enq_v,
        fifo6$in$enq__RDY,
        fifo6$out$first,
        fifo6$out$first__RDY);
    wire fifo7$out$deq__RDY;
    wire fifo7$in$enq__ENA;
    wire [95:0]fifo7$in$enq_v;
    wire fifo7$in$enq__RDY;
    wire [95:0]fifo7$out$first;
    wire fifo7$out$first__RDY;
    l_module_OC_FifoPong fifo7 (
        CLK,
        nRST,
        respond7__ENA_internal,
        fifo7$out$deq__RDY,
        fifo7$in$enq__ENA,
        fifo7$in$enq_v,
        fifo7$in$enq__RDY,
        fifo7$out$first,
        fifo7$out$first__RDY);
    wire fifo8$out$deq__RDY;
    wire fifo8$in$enq__ENA;
    wire [95:0]fifo8$in$enq_v;
    wire fifo8$in$enq__RDY;
    wire [95:0]fifo8$out$first;
    wire fifo8$out$first__RDY;
    l_module_OC_FifoPong fifo8 (
        CLK,
        nRST,
        respond8__ENA_internal,
        fifo8$out$deq__RDY,
        fifo8$in$enq__ENA,
        fifo8$in$enq_v,
        fifo8$in$enq__RDY,
        fifo8$out$first,
        fifo8$out$first__RDY);
    wire fifo9$out$deq__RDY;
    wire fifo9$in$enq__ENA;
    wire [95:0]fifo9$in$enq_v;
    wire fifo9$in$enq__RDY;
    wire [95:0]fifo9$out$first;
    wire fifo9$out$first__RDY;
    l_module_OC_FifoPong fifo9 (
        CLK,
        nRST,
        respond9__ENA_internal,
        fifo9$out$deq__RDY,
        fifo9$in$enq__ENA,
        fifo9$in$enq_v,
        fifo9$in$enq__RDY,
        fifo9$out$first,
        fifo9$out$first__RDY);
    wire fifo10$out$deq__ENA;
    wire fifo10$out$deq__RDY;
    wire fifo10$in$enq__ENA;
    wire [95:0]fifo10$in$enq_v;
    wire fifo10$in$enq__RDY;
    wire [95:0]fifo10$out$first;
    wire fifo10$out$first__RDY;
    l_module_OC_FifoPong fifo10 (
        CLK,
        nRST,
        fifo10$out$deq__ENA,
        fifo10$out$deq__RDY,
        fifo10$in$enq__ENA,
        fifo10$in$enq_v,
        fifo10$in$enq__RDY,
        fifo10$out$first,
        fifo10$out$first__RDY);
    reg[31:0] vsize;
    assign (in$say_meth == 0 ? &fifo0:in$say_meth == 1 ? &fifo1:in$say_meth == 2 ? &fifo2:in$say_meth == 3 ? &fifo3:in$say_meth == 4 ? &fifo4:in$say_meth == 5 ? &fifo5:in$say_meth == 6 ? &fifo6:in$say_meth == 7 ? &fifo7:in$say_meth == 8 ? &fifo8:&fifo9)$in$enq__ENA = in$say__ENA_internal;
    assign (in$say_meth == 0 ? &fifo0:in$say_meth == 1 ? &fifo1:in$say_meth == 2 ? &fifo2:in$say_meth == 3 ? &fifo3:in$say_meth == 4 ? &fifo4:in$say_meth == 5 ? &fifo5:in$say_meth == 6 ? &fifo6:in$say_meth == 7 ? &fifo7:in$say_meth == 8 ? &fifo8:&fifo9)$in$enq_v = temp;
    assign in$say__RDY = in$say__RDY_internal;
    assign in$say__RDY_internal = ((((((((fifo0$in$enq__RDY & fifo1$in$enq__RDY) & fifo2$in$enq__RDY) & fifo3$in$enq__RDY) & fifo4$in$enq__RDY) & fifo5$in$enq__RDY) & fifo6$in$enq__RDY) & fifo7$in$enq__RDY) & fifo8$in$enq__RDY) & fifo9$in$enq__RDY;
    assign ind$heard__ENA = respond0__ENA_internal || respond1__ENA_internal || respond2__ENA_internal || respond3__ENA_internal || respond4__ENA_internal || respond5__ENA_internal || respond6__ENA_internal || respond7__ENA_internal || respond8__ENA_internal || respond9__ENA_internal;
    assign ind$heard_heard_meth = respond0__ENA_internal ? 0 : respond1__ENA_internal ? 1 : respond2__ENA_internal ? 2 : respond3__ENA_internal ? 3 : respond4__ENA_internal ? 4 : respond5__ENA_internal ? 5 : respond6__ENA_internal ? 6 : respond7__ENA_internal ? 7 : respond8__ENA_internal ? 8 : 9;
    assign ind$heard_heard_v = respond0__ENA_internal ? temp$b : respond1__ENA_internal ? temp$b : respond2__ENA_internal ? temp$b : respond3__ENA_internal ? temp$b : respond4__ENA_internal ? temp$b : respond5__ENA_internal ? temp$b : respond6__ENA_internal ? temp$b : respond7__ENA_internal ? temp$b : respond8__ENA_internal ? temp$b : temp$b;
    assign respond0__RDY_internal = (fifo0$out$first__RDY & fifo0$out$deq__RDY) & ind$heard__RDY;
    assign respond1__RDY_internal = (fifo1$out$first__RDY & fifo1$out$deq__RDY) & ind$heard__RDY;
    assign respond2__RDY_internal = (fifo2$out$first__RDY & fifo2$out$deq__RDY) & ind$heard__RDY;
    assign respond3__RDY_internal = (fifo3$out$first__RDY & fifo3$out$deq__RDY) & ind$heard__RDY;
    assign respond4__RDY_internal = (fifo4$out$first__RDY & fifo4$out$deq__RDY) & ind$heard__RDY;
    assign respond5__RDY_internal = (fifo5$out$first__RDY & fifo5$out$deq__RDY) & ind$heard__RDY;
    assign respond6__RDY_internal = (fifo6$out$first__RDY & fifo6$out$deq__RDY) & ind$heard__RDY;
    assign respond7__RDY_internal = (fifo7$out$first__RDY & fifo7$out$deq__RDY) & ind$heard__RDY;
    assign respond8__RDY_internal = (fifo8$out$first__RDY & fifo8$out$deq__RDY) & ind$heard__RDY;
    assign respond9__RDY_internal = (fifo9$out$first__RDY & fifo9$out$deq__RDY) & ind$heard__RDY;
    assign temp$a = fifo9$out$first.a;
    assign temp$b = in$say_v;
    assign temp$c = fifo9$out$first.c;

    always @( posedge CLK) begin
      if (!nRST) begin
        vsize <= 0;
      end // nRST
    end // always @ (posedge CLK)
endmodule 

