`include "zynqTop.generated.vh"

`default_nettype none
module ZynqTop (
    output wire MAXIGP0_O$AR__ENA,
    output wire [31:0]MAXIGP0_O$AR$addr,
    output wire [11:0]MAXIGP0_O$AR$id,
    output wire [3:0]MAXIGP0_O$AR$len,
    input wire MAXIGP0_O$AR__RDY,
    output wire MAXIGP0_O$AW__ENA,
    output wire [31:0]MAXIGP0_O$AW$addr,
    output wire [11:0]MAXIGP0_O$AW$id,
    output wire [3:0]MAXIGP0_O$AW$len,
    input wire MAXIGP0_O$AW__RDY,
    output wire MAXIGP0_O$W__ENA,
    output wire [31:0]MAXIGP0_O$W$data,
    output wire [11:0]MAXIGP0_O$W$id,
    output wire MAXIGP0_O$W$last,
    input wire MAXIGP0_O$W__RDY,
    input wire MAXIGP0_I$B__ENA,
    input wire [11:0]MAXIGP0_I$B$id,
    input wire [1:0]MAXIGP0_I$B$resp,
    output wire MAXIGP0_I$B__RDY,
    input wire MAXIGP0_I$R__ENA,
    input wire [31:0]MAXIGP0_I$R$data,
    input wire [11:0]MAXIGP0_I$R$id,
    input wire MAXIGP0_I$R$last,
    input wire [1:0]MAXIGP0_I$R$resp,
    output wire MAXIGP0_I$R__RDY,
    input wire CLK,
    input wire nRST,
    inout wire [14:0]DDR_Addr,
    inout wire [2:0]DDR_BankAddr,
    inout wire DDR_CAS_n,
    inout wire DDR_CKE,
    inout wire DDR_Clk_n,
    inout wire DDR_Clk_p,
    inout wire DDR_CS_n,
    inout wire [3:0]DDR_DM,
    inout wire [31:0]DDR_DQ,
    inout wire [3:0]DDR_DQS_n,
    inout wire [3:0]DDR_DQS_p,
    inout wire DDR_DRSTB,
    inout wire DDR_ODT,
    inout wire DDR_RAS_n,
    inout wire FIXED_IO_ddr_vrn,
    inout wire FIXED_IO_ddr_vrp,
    inout wire DDR_WEB,
    inout wire FIXED_IO_ps_clk,
    inout wire FIXED_IO_ps_porb,
    inout wire FIXED_IO_ps_srstb,
    input wire interrupt,
    inout wire [53:0]MIO,
    output wire [3:0]FCLKCLK,
    input wire [3:0]FCLKCLKTRIGN,
    output wire [3:0]FCLKRESETN);
    wire RULEinit__ENA;
    assign RULEinit__ENA = 1;
    P7Wrap zt (
        .MAXIGP0_O$AR__ENA(MAXIGP0_O$AR__ENA),
        .MAXIGP0_O$AR$addr(MAXIGP0_O$AR$addr),
        .MAXIGP0_O$AR$id(MAXIGP0_O$AR$id),
        .MAXIGP0_O$AR$len(MAXIGP0_O$AR$len),
        .MAXIGP0_O$AR__RDY(MAXIGP0_O$AR__RDY),
        .MAXIGP0_O$AW__ENA(MAXIGP0_O$AW__ENA),
        .MAXIGP0_O$AW$addr(MAXIGP0_O$AW$addr),
        .MAXIGP0_O$AW$id(MAXIGP0_O$AW$id),
        .MAXIGP0_O$AW$len(MAXIGP0_O$AW$len),
        .MAXIGP0_O$AW__RDY(MAXIGP0_O$AW__RDY),
        .MAXIGP0_O$W__ENA(MAXIGP0_O$W__ENA),
        .MAXIGP0_O$W$data(MAXIGP0_O$W$data),
        .MAXIGP0_O$W$id(MAXIGP0_O$W$id),
        .MAXIGP0_O$W$last(MAXIGP0_O$W$last),
        .MAXIGP0_O$W__RDY(MAXIGP0_O$W__RDY),
        .MAXIGP0_I$B__ENA(MAXIGP0_I$B__ENA),
        .MAXIGP0_I$B$id(MAXIGP0_I$B$id),
        .MAXIGP0_I$B$resp(MAXIGP0_I$B$resp),
        .MAXIGP0_I$B__RDY(MAXIGP0_I$B__RDY),
        .MAXIGP0_I$R__ENA(MAXIGP0_I$R__ENA),
        .MAXIGP0_I$R$data(MAXIGP0_I$R$data),
        .MAXIGP0_I$R$id(MAXIGP0_I$R$id),
        .MAXIGP0_I$R$last(MAXIGP0_I$R$last),
        .MAXIGP0_I$R$resp(MAXIGP0_I$R$resp),
        .MAXIGP0_I$R__RDY(MAXIGP0_I$R__RDY),
        .CLK(CLK),
        .nRST(nRST),
        .DDR_Addr(DDR_Addr),
        .DDR_BankAddr(DDR_BankAddr),
        .DDR_CAS_n(DDR_CAS_n),
        .DDR_CKE(DDR_CKE),
        .DDR_Clk_n(DDR_Clk_n),
        .DDR_Clk_p(DDR_Clk_p),
        .DDR_CS_n(DDR_CS_n),
        .DDR_DM(DDR_DM),
        .DDR_DQ(DDR_DQ),
        .DDR_DQS_n(DDR_DQS_n),
        .DDR_DQS_p(DDR_DQS_p),
        .DDR_DRSTB(DDR_DRSTB),
        .DDR_ODT(DDR_ODT),
        .DDR_RAS_n(DDR_RAS_n),
        .FIXED_IO_ddr_vrn(FIXED_IO_ddr_vrn),
        .FIXED_IO_ddr_vrp(FIXED_IO_ddr_vrp),
        .DDR_WEB(DDR_WEB),
        .FIXED_IO_ps_clk(FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb(FIXED_IO_ps_porb),
        .FIXED_IO_ps_srstb(FIXED_IO_ps_srstb),
        .interrupt(interrupt),
        .MIO(MIO),
        .FCLKCLK(FCLKCLK),
        .FCLKCLKTRIGN(FCLKCLKTRIGN),
        .FCLKRESETN(FCLKRESETN));
endmodule 

`default_nettype wire    // set back to default value
