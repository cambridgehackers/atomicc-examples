`ifndef __grayCounter_GENERATED__VH__
`define __grayCounter_GENERATED__VH__

//METASTART; GrayCounter
//METAGUARD; increment; 1;
//METAGUARD; decrement; 1;
//METAGUARD; readGray; 1;
//METAGUARD; writeGray; 1;
//METAGUARD; readBin; 1;
//METAGUARD; writeBin; 1;
//METAGUARD; RULE$incdec; increment__ENA != decrement__ENA;
//METAGUARD; RULE$init; 1;
//METARULES; RULE$incdec; RULE$init
`endif
