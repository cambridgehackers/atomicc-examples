`ifndef __gearNto1_GENERATED__VH__
`define __gearNto1_GENERATED__VH__

//METASTART; GearNto1Base
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; ( !( 0 == ( ( c != 0 ) ^ 1 ) ) );
//METAGUARD; out$deq; ( !( 0 == ( ( c == 0 ) ^ 1 ) ) );
//METAGUARD; out$first; ( !( 0 == ( ( c == 0 ) ^ 1 ) ) );
`endif
