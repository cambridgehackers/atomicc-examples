`ifndef __axiTop_GENERATED__VH__
`define __axiTop_GENERATED__VH__

//METASTART; AxiTop
//METAINTERNAL; reqArs; Fifo1Base(width=6);
//METAINTERNAL; reqAws; Fifo1Base(width=6);
//METAINTERNAL; writeDone; Fifo1Base(width=6);
//METAINTERNAL; requestValue; Fifo1Base(width=32);
//METAINTERNAL; readData; Fifo1Base(width=38);
//METAINTERNAL; writeData; Fifo1Base(width=32);
//METAINTERNAL; user; UserTop;
//METAINVOKE; MAXIGP0_O$AR__ENA; :reqArs$in$enq__ENA;
//METAEXCLUSIVE; MAXIGP0_O$AR__ENA; RULE$lread__ENA
//METAGUARD; MAXIGP0_O$AR; reqArs$in$enq__RDY;
//METAINVOKE; MAXIGP0_O$AW__ENA; :reqAws$in$enq__ENA;
//METAEXCLUSIVE; MAXIGP0_O$AW__ENA; RULE$lwrite__ENA
//METAGUARD; MAXIGP0_O$AW; reqAws$in$enq__RDY;
//METAINVOKE; MAXIGP0_O$W__ENA; :writeData$in$enq__ENA;
//METAGUARD; MAXIGP0_O$W; writeData$in$enq__RDY;
//METAINVOKE; readUser$enq__ENA; :requestValue$in$enq__ENA;
//METAGUARD; readUser$enq; requestValue$in$enq__RDY;
//METABEFORE; RULE$init__ENA; :RULE$lwrite__ENA
//METAGUARD; RULE$init; 1;
//METAINVOKE; RULE$lread__ENA; 1:readData$in$enq__ENA;readCount == 0:reqArs$out$deq__ENA;:reqArs$out$first;!( portalRControl || ( !( readAddr == 0 ) ) ):requestValue$out$deq__ENA;!( portalRControl || ( !( readAddr == 0 ) ) ):requestValue$out$first;
//METABEFORE; RULE$lread__ENA; :MAXIGP0_O$AR__ENA
//METAGUARD; RULE$lread; reqArs$out$first__RDY && ( ( portalRControl && readData$in$enq__RDY && ( reqArs$out$deq__RDY || ( !( readCount == 0 ) ) ) ) || ( ( !portalRControl ) && readData$in$enq__RDY && ( ( requestValue$out$first__RDY && ( ( requestValue$out$deq__RDY && ( reqArs$out$deq__RDY || ( !( readCount == 0 ) ) ) ) || ( ( !requestValue$out$deq__RDY ) && ( !( ( readAddr == 0 ) || ( !( reqArs$out$deq__RDY || ( !( readCount == 0 ) ) ) ) ) ) ) ) ) || ( ( !requestValue$out$first__RDY ) && ( !( ( readAddr == 0 ) || ( !( reqArs$out$deq__RDY || ( !( readCount == 0 ) ) ) ) ) ) ) ) ) );
//METAINVOKE; RULE$lreadData__ENA; :MAXIGP0_I$R__ENA;:readData$out$deq__ENA;:readData$out$first;
//METAGUARD; RULE$lreadData; readData$out$first__RDY && MAXIGP0_I$R__RDY && readData$out$deq__RDY;
//METAINVOKE; RULE$lwrite__ENA; writeCount == 0:reqAws$out$deq__ENA;:reqAws$out$first;!portalWControl:user$write$enq__ENA;:writeData$out$deq__ENA;:writeData$out$first;writeCount == 0:writeDone$in$enq__ENA;
//METABEFORE; RULE$lwrite__ENA; :MAXIGP0_O$AW__ENA
//METAGUARD; RULE$lwrite; reqAws$out$first__RDY && writeData$out$first__RDY && ( ( portalWControl && writeData$out$deq__RDY && ( ( writeDone$in$enq__RDY && ( reqAws$out$deq__RDY || ( !( writeCount == 0 ) ) ) ) || ( ( !writeDone$in$enq__RDY ) && ( !( writeCount == 0 ) ) ) ) ) || ( ( !portalWControl ) && writeData$out$deq__RDY && ( ( writeDone$in$enq__RDY && ( ( ( writeCount == 0 ) && user$write$enq__RDY && reqAws$out$deq__RDY ) || ( ( !( writeCount == 0 ) ) && user$write$enq__RDY ) ) ) || ( ( !writeDone$in$enq__RDY ) && ( !( ( writeCount == 0 ) || ( !user$write$enq__RDY ) ) ) ) ) ) );
//METAINVOKE; RULE$writeResponse__ENA; :MAXIGP0_I$B__ENA;:writeDone$out$deq__ENA;:writeDone$out$first;
//METAGUARD; RULE$writeResponse; writeDone$out$first__RDY && MAXIGP0_I$B__RDY && writeDone$out$deq__RDY;
//METARULES; RULE$init; RULE$lread; RULE$lreadData; RULE$lwrite; RULE$writeResponse
//METACONNECT; readUser$enq__ENA; user$read$enq__ENA
//METACONNECT; readUser$enq__RDY; user$read$enq__RDY
`endif
