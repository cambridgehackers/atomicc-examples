
    assign bscan$toBscan.enq$v = test.__traceMemory$out.first;
    assign bscan$toBscan.enq__ENA = test.__traceMemory$out.first__RDY;
    assign test.__traceMemory$out.deq__ENA = readUser.enq__ENA;
