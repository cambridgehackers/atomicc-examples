`ifndef __syncFF_GENERATED__VH__
`define __syncFF_GENERATED__VH__

//METASTART; SyncFF
//METAGUARD; RULE$init; 1;
//METARULES; RULE$init
`endif
