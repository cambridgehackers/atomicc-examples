`include "atomicclib.vh"

//METASTART; ResetInverter
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$init
