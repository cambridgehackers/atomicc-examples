`ifndef __resetInverter_GENERATED__VH__
`define __resetInverter_GENERATED__VH__

//METASTART; ResetInverter
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$init
`endif
