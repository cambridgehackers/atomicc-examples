`include "atomicc.generated.vh"
`default_nettype none
module P7Wrap (
    inout wire [54 - 1:0]MIO,
    inout wire [15 - 1:0]DDR_Addr,
    inout wire [3 - 1:0]DDR_BankAddr,
    inout wire DDR_CAS_n,
    inout wire DDR_CKE,
    inout wire DDR_Clk_n,
    inout wire DDR_Clk_p,
    inout wire DDR_CS_n,
    inout wire [4 - 1:0]DDR_DM,
    inout wire [32 - 1:0]DDR_DQ,
    inout wire [4 - 1:0]DDR_DQS_n,
    inout wire [4 - 1:0]DDR_DQS_p,
    inout wire DDR_DRSTB,
    inout wire DDR_ODT,
    inout wire DDR_RAS_n,
    inout wire FIXED_IO_ddr_vrn,
    inout wire FIXED_IO_ddr_vrp,
    inout wire DDR_WEB,
    inout wire FIXED_IO_ps_clk,
    inout wire FIXED_IO_ps_porb,
    inout wire FIXED_IO_ps_srstb,
    ZynqInterrupt.server intr,
    MaxiO.client MAXIGP0_O,
    MaxiI.server MAXIGP0_I,
    Pps7fclk.server FCLK,
    inout wire i2c0$scl,
    inout wire i2c0$sda,
    inout wire i2c1$scl,
    inout wire i2c1$sda);
    logic CLK;
    logic nRST;
    logic pps$EMIOI2C0SCLO;
    logic pps$EMIOI2C0SCLTN;
    logic pps$EMIOI2C0SDAO;
    logic pps$EMIOI2C0SDATN;
    logic pps$EMIOI2C1SCLO;
    logic pps$EMIOI2C1SCLTN;
    logic pps$EMIOI2C1SDAO;
    logic pps$EMIOI2C1SDATN;
    logic pps$MAXIGP0WLAST;
    logic tscl0$O;
    logic tscl1$O;
    logic tsda0$O;
    logic tsda1$O;
    PS7 pps (
        .MIO(MIO),
        .DDRA(DDR_Addr),
        .DDRARB(4'd0),
        .DDRBA(DDR_BankAddr),
        .DDRCASB(DDR_CAS_n),
        .DDRCKE(DDR_CKE),
        .DDRCKN(DDR_Clk_n),
        .DDRCKP(DDR_Clk_p),
        .DDRCSB(DDR_CS_n),
        .DDRDM(DDR_DM),
        .DDRDQ(DDR_DQ),
        .DDRDQSN(DDR_DQS_n),
        .DDRDQSP(DDR_DQS_p),
        .DDRDRSTB(DDR_DRSTB),
        .DDRODT(DDR_ODT),
        .DDRRASB(DDR_RAS_n),
        .DDRVRN(FIXED_IO_ddr_vrn),
        .DDRVRP(FIXED_IO_ddr_vrp),
        .DDRWEB(DDR_WEB),
        .DMA0ACLK(1'd0),
        .DMA0DAREADY(1'd0),
        .DMA0DATYPE(),
        .DMA0DAVALID(),
        .DMA0DRLAST(1'd0),
        .DMA0DRREADY(),
        .DMA0DRTYPE(2'd0),
        .DMA0DRVALID(1'd0),
        .DMA0RSTN(),
        .DMA1ACLK(1'd0),
        .DMA1DAREADY(1'd0),
        .DMA1DATYPE(),
        .DMA1DAVALID(),
        .DMA1DRLAST(1'd0),
        .DMA1DRREADY(),
        .DMA1DRTYPE(2'd0),
        .DMA1DRVALID(1'd0),
        .DMA1RSTN(),
        .DMA2ACLK(1'd0),
        .DMA2DAREADY(1'd0),
        .DMA2DATYPE(),
        .DMA2DAVALID(),
        .DMA2DRLAST(1'd0),
        .DMA2DRREADY(),
        .DMA2DRTYPE(2'd0),
        .DMA2DRVALID(1'd0),
        .DMA2RSTN(),
        .DMA3ACLK(1'd0),
        .DMA3DAREADY(1'd0),
        .DMA3DATYPE(),
        .DMA3DAVALID(),
        .DMA3DRLAST(1'd0),
        .DMA3DRREADY(),
        .DMA3DRTYPE(2'd0),
        .DMA3DRVALID(1'd0),
        .DMA3RSTN(),
        .EMIOCAN0PHYRX(1'd0),
        .EMIOCAN0PHYTX(),
        .EMIOCAN1PHYRX(1'd0),
        .EMIOCAN1PHYTX(),
        .EMIOENET0EXTINTIN(1'd0),
        .EMIOENET0GMIICOL(1'd0),
        .EMIOENET0GMIICRS(1'd0),
        .EMIOENET0GMIIRXCLK(1'd0),
        .EMIOENET0GMIIRXD(8'd0),
        .EMIOENET0GMIIRXDV(1'd0),
        .EMIOENET0GMIIRXER(1'd0),
        .EMIOENET0GMIITXCLK(1'd0),
        .EMIOENET0GMIITXD(),
        .EMIOENET0GMIITXEN(),
        .EMIOENET0GMIITXER(),
        .EMIOENET0MDIOI(1'd0),
        .EMIOENET0MDIOMDC(),
        .EMIOENET0MDIOO(),
        .EMIOENET0MDIOTN(),
        .EMIOENET0PTPDELAYREQRX(),
        .EMIOENET0PTPDELAYREQTX(),
        .EMIOENET0PTPPDELAYREQRX(),
        .EMIOENET0PTPPDELAYREQTX(),
        .EMIOENET0PTPPDELAYRESPRX(),
        .EMIOENET0PTPPDELAYRESPTX(),
        .EMIOENET0PTPSYNCFRAMERX(),
        .EMIOENET0PTPSYNCFRAMETX(),
        .EMIOENET0SOFRX(),
        .EMIOENET0SOFTX(),
        .EMIOENET1EXTINTIN(1'd0),
        .EMIOENET1GMIICOL(1'd0),
        .EMIOENET1GMIICRS(1'd0),
        .EMIOENET1GMIIRXCLK(1'd0),
        .EMIOENET1GMIIRXD(8'd0),
        .EMIOENET1GMIIRXDV(1'd0),
        .EMIOENET1GMIIRXER(1'd0),
        .EMIOENET1GMIITXCLK(1'd0),
        .EMIOENET1GMIITXD(),
        .EMIOENET1GMIITXEN(),
        .EMIOENET1GMIITXER(),
        .EMIOENET1MDIOI(1'd0),
        .EMIOENET1MDIOMDC(),
        .EMIOENET1MDIOO(),
        .EMIOENET1MDIOTN(),
        .EMIOENET1PTPDELAYREQRX(),
        .EMIOENET1PTPDELAYREQTX(),
        .EMIOENET1PTPPDELAYREQRX(),
        .EMIOENET1PTPPDELAYREQTX(),
        .EMIOENET1PTPPDELAYRESPRX(),
        .EMIOENET1PTPPDELAYRESPTX(),
        .EMIOENET1PTPSYNCFRAMERX(),
        .EMIOENET1PTPSYNCFRAMETX(),
        .EMIOENET1SOFRX(),
        .EMIOENET1SOFTX(),
        .EMIOGPIOI(64'd0),
        .EMIOGPIOO(),
        .EMIOGPIOTN(),
        .EMIOI2C0SCLI(tscl0$O),
        .EMIOI2C0SCLO(pps$EMIOI2C0SCLO),
        .EMIOI2C0SCLTN(pps$EMIOI2C0SCLTN),
        .EMIOI2C0SDAI(tsda0$O),
        .EMIOI2C0SDAO(pps$EMIOI2C0SDAO),
        .EMIOI2C0SDATN(pps$EMIOI2C0SDATN),
        .EMIOI2C1SCLI(tscl1$O),
        .EMIOI2C1SCLO(pps$EMIOI2C1SCLO),
        .EMIOI2C1SCLTN(pps$EMIOI2C1SCLTN),
        .EMIOI2C1SDAI(tsda1$O),
        .EMIOI2C1SDAO(pps$EMIOI2C1SDAO),
        .EMIOI2C1SDATN(pps$EMIOI2C1SDATN),
        .EMIOPJTAGTCK(1'd0),
        .EMIOPJTAGTDI(1'd0),
        .EMIOPJTAGTDO(),
        .EMIOPJTAGTDTN(),
        .EMIOPJTAGTMS(1'd0),
        .EMIOSDIO0BUSPOW(),
        .EMIOSDIO0BUSVOLT(),
        .EMIOSDIO0CDN(1'd0),
        .EMIOSDIO0CLK(),
        .EMIOSDIO0CLKFB(1'd0),
        .EMIOSDIO0CMDI(1'd0),
        .EMIOSDIO0CMDO(),
        .EMIOSDIO0CMDTN(),
        .EMIOSDIO0DATAI(4'd0),
        .EMIOSDIO0DATAO(),
        .EMIOSDIO0DATATN(),
        .EMIOSDIO0LED(),
        .EMIOSDIO0WP(1'd0),
        .EMIOSDIO1BUSPOW(),
        .EMIOSDIO1BUSVOLT(),
        .EMIOSDIO1CDN(1'd0),
        .EMIOSDIO1CLK(),
        .EMIOSDIO1CLKFB(1'd0),
        .EMIOSDIO1CMDI(1'd0),
        .EMIOSDIO1CMDO(),
        .EMIOSDIO1CMDTN(),
        .EMIOSDIO1DATAI(4'd0),
        .EMIOSDIO1DATAO(),
        .EMIOSDIO1DATATN(),
        .EMIOSDIO1LED(),
        .EMIOSDIO1WP(1'd0),
        .EMIOSPI0MI(1'd0),
        .EMIOSPI0MO(),
        .EMIOSPI0MOTN(),
        .EMIOSPI0SCLKI(1'd0),
        .EMIOSPI0SCLKO(),
        .EMIOSPI0SCLKTN(),
        .EMIOSPI0SI(1'd0),
        .EMIOSPI0SO(),
        .EMIOSPI0SSIN(1'd0),
        .EMIOSPI0SSNTN(),
        .EMIOSPI0SSON(),
        .EMIOSPI0STN(),
        .EMIOSPI1MI(1'd0),
        .EMIOSPI1MO(),
        .EMIOSPI1MOTN(),
        .EMIOSPI1SCLKI(1'd0),
        .EMIOSPI1SCLKO(),
        .EMIOSPI1SCLKTN(),
        .EMIOSPI1SI(1'd0),
        .EMIOSPI1SO(),
        .EMIOSPI1SSIN(1'd0),
        .EMIOSPI1SSNTN(),
        .EMIOSPI1SSON(),
        .EMIOSPI1STN(),
        .EMIOSRAMINTIN(1'd0),
        .EMIOTRACECLK(1'd0),
        .EMIOTRACECTL(),
        .EMIOTRACEDATA(),
        .EMIOTTC0CLKI(3'd0),
        .EMIOTTC0WAVEO(),
        .EMIOTTC1CLKI(3'd0),
        .EMIOTTC1WAVEO(),
        .EMIOUART0CTSN(1'd0),
        .EMIOUART0DCDN(1'd0),
        .EMIOUART0DSRN(1'd0),
        .EMIOUART0DTRN(),
        .EMIOUART0RIN(1'd0),
        .EMIOUART0RTSN(),
        .EMIOUART0RX(1'd0),
        .EMIOUART0TX(),
        .EMIOUART1CTSN(1'd0),
        .EMIOUART1DCDN(1'd0),
        .EMIOUART1DSRN(1'd0),
        .EMIOUART1DTRN(),
        .EMIOUART1RIN(1'd0),
        .EMIOUART1RTSN(),
        .EMIOUART1RX(1'd0),
        .EMIOUART1TX(),
        .EMIOUSB0PORTINDCTL(),
        .EMIOUSB0VBUSPWRFAULT(1'd0),
        .EMIOUSB0VBUSPWRSELECT(),
        .EMIOUSB1PORTINDCTL(),
        .EMIOUSB1VBUSPWRFAULT(1'd0),
        .EMIOUSB1VBUSPWRSELECT(),
        .EMIOWDTCLKI(1'd0),
        .EMIOWDTRSTO(),
        .EVENTEVENTI(1'd0),
        .EVENTEVENTO(),
        .EVENTSTANDBYWFE(),
        .EVENTSTANDBYWFI(),
        .FCLKCLK(FCLK.CLK),
        .FCLKCLKTRIGN(FCLK.CLKTRIGN),
        .FCLKRESETN(FCLK.RESETN),
        .FPGAIDLEN(1'd1),
        .FTMDTRACEINATID(4'd0),
        .FTMDTRACEINCLOCK(1'd0),
        .FTMDTRACEINDATA(32'd0),
        .FTMDTRACEINVALID(1'd0),
        .FTMTF2PDEBUG(32'd0),
        .FTMTF2PTRIG(4'd0),
        .FTMTF2PTRIGACK(),
        .FTMTP2FDEBUG(),
        .FTMTP2FTRIG(),
        .FTMTP2FTRIGACK(4'd0),
        .IRQF2P(intr.interrupt),
        .IRQP2F(),
        .MAXIGP0ACLK(CLK),
        .MAXIGP0ARADDR(MAXIGP0_O.AR$addr),
        .MAXIGP0ARBURST(),
        .MAXIGP0ARCACHE(),
        .MAXIGP0ARESETN(),
        .MAXIGP0ARID(MAXIGP0_O.AR$id),
        .MAXIGP0ARLEN(MAXIGP0_O.AR$len),
        .MAXIGP0ARLOCK(),
        .MAXIGP0ARPROT(),
        .MAXIGP0ARQOS(),
        .MAXIGP0ARREADY(MAXIGP0_O.AR__RDY),
        .MAXIGP0ARSIZE(),
        .MAXIGP0ARVALID(MAXIGP0_O.AR__ENA),
        .MAXIGP0AWADDR(MAXIGP0_O.AW$addr),
        .MAXIGP0AWBURST(),
        .MAXIGP0AWCACHE(),
        .MAXIGP0AWID(MAXIGP0_O.AW$id),
        .MAXIGP0AWLEN(MAXIGP0_O.AW$len),
        .MAXIGP0AWLOCK(),
        .MAXIGP0AWPROT(),
        .MAXIGP0AWQOS(),
        .MAXIGP0AWREADY(MAXIGP0_O.AW__RDY),
        .MAXIGP0AWSIZE(),
        .MAXIGP0AWVALID(MAXIGP0_O.AW__ENA),
        .MAXIGP0BID(MAXIGP0_I.B__ENA ? MAXIGP0_I.B$id : 12'd0),
        .MAXIGP0BREADY(MAXIGP0_I.B__RDY),
        .MAXIGP0BRESP(MAXIGP0_I.B__ENA ? MAXIGP0_I.B$resp : 2'd0),
        .MAXIGP0BVALID(MAXIGP0_I.B__ENA),
        .MAXIGP0RDATA(MAXIGP0_I.R__ENA ? MAXIGP0_I.R$data : 32'd0),
        .MAXIGP0RID(MAXIGP0_I.R__ENA ? MAXIGP0_I.R$id : 12'd0),
        .MAXIGP0RLAST(MAXIGP0_I.R__ENA && MAXIGP0_I.R$last),
        .MAXIGP0RREADY(MAXIGP0_I.R__RDY),
        .MAXIGP0RRESP(MAXIGP0_I.R__ENA ? MAXIGP0_I.R$resp : 2'd0),
        .MAXIGP0RVALID(MAXIGP0_I.R__ENA),
        .MAXIGP0WDATA(MAXIGP0_O.W$data),
        .MAXIGP0WID(MAXIGP0_O.W$id),
        .MAXIGP0WLAST(pps$MAXIGP0WLAST),
        .MAXIGP0WREADY(MAXIGP0_O.W__RDY),
        .MAXIGP0WSTRB(),
        .MAXIGP0WVALID(MAXIGP0_O.W__ENA),
        .MAXIGP1ACLK(1'd0),
        .MAXIGP1ARADDR(),
        .MAXIGP1ARBURST(),
        .MAXIGP1ARCACHE(),
        .MAXIGP1ARESETN(),
        .MAXIGP1ARID(),
        .MAXIGP1ARLEN(),
        .MAXIGP1ARLOCK(),
        .MAXIGP1ARPROT(),
        .MAXIGP1ARQOS(),
        .MAXIGP1ARREADY(1'd0),
        .MAXIGP1ARSIZE(),
        .MAXIGP1ARVALID(),
        .MAXIGP1AWADDR(),
        .MAXIGP1AWBURST(),
        .MAXIGP1AWCACHE(),
        .MAXIGP1AWID(),
        .MAXIGP1AWLEN(),
        .MAXIGP1AWLOCK(),
        .MAXIGP1AWPROT(),
        .MAXIGP1AWQOS(),
        .MAXIGP1AWREADY(1'd0),
        .MAXIGP1AWSIZE(),
        .MAXIGP1AWVALID(),
        .MAXIGP1BID(12'd0),
        .MAXIGP1BREADY(),
        .MAXIGP1BRESP(2'd0),
        .MAXIGP1BVALID(1'd0),
        .MAXIGP1RDATA(32'd0),
        .MAXIGP1RID(12'd0),
        .MAXIGP1RLAST(1'd0),
        .MAXIGP1RREADY(),
        .MAXIGP1RRESP(2'd0),
        .MAXIGP1RVALID(1'd0),
        .MAXIGP1WDATA(),
        .MAXIGP1WID(),
        .MAXIGP1WLAST(),
        .MAXIGP1WREADY(1'd0),
        .MAXIGP1WSTRB(),
        .MAXIGP1WVALID(),
        .PSCLK(FIXED_IO_ps_clk),
        .PSPORB(FIXED_IO_ps_porb),
        .PSSRSTB(FIXED_IO_ps_srstb),
        .SAXIACPACLK(1'd0),
        .SAXIACPARADDR(32'd0),
        .SAXIACPARBURST(2'd0),
        .SAXIACPARCACHE(4'd0),
        .SAXIACPARESETN(),
        .SAXIACPARID(3'd0),
        .SAXIACPARLEN(4'd0),
        .SAXIACPARLOCK(2'd0),
        .SAXIACPARPROT(3'd0),
        .SAXIACPARQOS(4'd0),
        .SAXIACPARREADY(),
        .SAXIACPARSIZE(2'd0),
        .SAXIACPARUSER(5'd0),
        .SAXIACPARVALID(1'd0),
        .SAXIACPAWADDR(32'd0),
        .SAXIACPAWBURST(2'd0),
        .SAXIACPAWCACHE(4'd0),
        .SAXIACPAWID(3'd0),
        .SAXIACPAWLEN(4'd0),
        .SAXIACPAWLOCK(2'd0),
        .SAXIACPAWPROT(3'd0),
        .SAXIACPAWQOS(4'd0),
        .SAXIACPAWREADY(),
        .SAXIACPAWSIZE(2'd0),
        .SAXIACPAWUSER(5'd0),
        .SAXIACPAWVALID(1'd0),
        .SAXIACPBID(),
        .SAXIACPBREADY(1'd0),
        .SAXIACPBRESP(),
        .SAXIACPBVALID(),
        .SAXIACPRDATA(),
        .SAXIACPRID(),
        .SAXIACPRLAST(),
        .SAXIACPRREADY(1'd0),
        .SAXIACPRRESP(),
        .SAXIACPRVALID(),
        .SAXIACPWDATA(64'd0),
        .SAXIACPWID(3'd0),
        .SAXIACPWLAST(1'd0),
        .SAXIACPWREADY(),
        .SAXIACPWSTRB(8'd0),
        .SAXIACPWVALID(1'd0),
        .SAXIGP0ACLK(1'd0),
        .SAXIGP0ARADDR(32'd0),
        .SAXIGP0ARBURST(2'd0),
        .SAXIGP0ARCACHE(4'd0),
        .SAXIGP0ARESETN(),
        .SAXIGP0ARID(6'd0),
        .SAXIGP0ARLEN(4'd0),
        .SAXIGP0ARLOCK(2'd0),
        .SAXIGP0ARPROT(3'd0),
        .SAXIGP0ARQOS(4'd0),
        .SAXIGP0ARREADY(),
        .SAXIGP0ARSIZE(2'd0),
        .SAXIGP0ARVALID(1'd0),
        .SAXIGP0AWADDR(32'd0),
        .SAXIGP0AWBURST(2'd0),
        .SAXIGP0AWCACHE(4'd0),
        .SAXIGP0AWID(6'd0),
        .SAXIGP0AWLEN(4'd0),
        .SAXIGP0AWLOCK(2'd0),
        .SAXIGP0AWPROT(3'd0),
        .SAXIGP0AWQOS(4'd0),
        .SAXIGP0AWREADY(),
        .SAXIGP0AWSIZE(2'd0),
        .SAXIGP0AWVALID(1'd0),
        .SAXIGP0BID(),
        .SAXIGP0BREADY(1'd0),
        .SAXIGP0BRESP(),
        .SAXIGP0BVALID(),
        .SAXIGP0RDATA(),
        .SAXIGP0RID(),
        .SAXIGP0RLAST(),
        .SAXIGP0RREADY(1'd0),
        .SAXIGP0RRESP(),
        .SAXIGP0RVALID(),
        .SAXIGP0WDATA(32'd0),
        .SAXIGP0WID(6'd0),
        .SAXIGP0WLAST(1'd0),
        .SAXIGP0WREADY(),
        .SAXIGP0WSTRB(4'd0),
        .SAXIGP0WVALID(1'd0),
        .SAXIGP1ACLK(1'd0),
        .SAXIGP1ARADDR(32'd0),
        .SAXIGP1ARBURST(2'd0),
        .SAXIGP1ARCACHE(4'd0),
        .SAXIGP1ARESETN(),
        .SAXIGP1ARID(6'd0),
        .SAXIGP1ARLEN(4'd0),
        .SAXIGP1ARLOCK(2'd0),
        .SAXIGP1ARPROT(3'd0),
        .SAXIGP1ARQOS(4'd0),
        .SAXIGP1ARREADY(),
        .SAXIGP1ARSIZE(2'd0),
        .SAXIGP1ARVALID(1'd0),
        .SAXIGP1AWADDR(32'd0),
        .SAXIGP1AWBURST(2'd0),
        .SAXIGP1AWCACHE(4'd0),
        .SAXIGP1AWID(6'd0),
        .SAXIGP1AWLEN(4'd0),
        .SAXIGP1AWLOCK(2'd0),
        .SAXIGP1AWPROT(3'd0),
        .SAXIGP1AWQOS(4'd0),
        .SAXIGP1AWREADY(),
        .SAXIGP1AWSIZE(2'd0),
        .SAXIGP1AWVALID(1'd0),
        .SAXIGP1BID(),
        .SAXIGP1BREADY(1'd0),
        .SAXIGP1BRESP(),
        .SAXIGP1BVALID(),
        .SAXIGP1RDATA(),
        .SAXIGP1RID(),
        .SAXIGP1RLAST(),
        .SAXIGP1RREADY(1'd0),
        .SAXIGP1RRESP(),
        .SAXIGP1RVALID(),
        .SAXIGP1WDATA(32'd0),
        .SAXIGP1WID(6'd0),
        .SAXIGP1WLAST(1'd0),
        .SAXIGP1WREADY(),
        .SAXIGP1WSTRB(4'd0),
        .SAXIGP1WVALID(1'd0),
        .SAXIHP0ACLK(1'd0),
        .SAXIHP0ARADDR(32'd0),
        .SAXIHP0ARBURST(2'd0),
        .SAXIHP0ARCACHE(4'd0),
        .SAXIHP0ARESETN(),
        .SAXIHP0ARID(6'd0),
        .SAXIHP0ARLEN(4'd0),
        .SAXIHP0ARLOCK(2'd0),
        .SAXIHP0ARPROT(3'd0),
        .SAXIHP0ARQOS(4'd0),
        .SAXIHP0ARREADY(),
        .SAXIHP0ARSIZE(2'd0),
        .SAXIHP0ARVALID(1'd0),
        .SAXIHP0AWADDR(32'd0),
        .SAXIHP0AWBURST(2'd0),
        .SAXIHP0AWCACHE(4'd0),
        .SAXIHP0AWID(6'd0),
        .SAXIHP0AWLEN(4'd0),
        .SAXIHP0AWLOCK(2'd0),
        .SAXIHP0AWPROT(3'd0),
        .SAXIHP0AWQOS(4'd0),
        .SAXIHP0AWREADY(),
        .SAXIHP0AWSIZE(2'd0),
        .SAXIHP0AWVALID(1'd0),
        .SAXIHP0BID(),
        .SAXIHP0BREADY(1'd0),
        .SAXIHP0BRESP(),
        .SAXIHP0BVALID(),
        .SAXIHP0RACOUNT(),
        .SAXIHP0RCOUNT(),
        .SAXIHP0RDATA(),
        .SAXIHP0RDISSUECAP1EN(1'd0),
        .SAXIHP0RID(),
        .SAXIHP0RLAST(),
        .SAXIHP0RREADY(1'd0),
        .SAXIHP0RRESP(),
        .SAXIHP0RVALID(),
        .SAXIHP0WACOUNT(),
        .SAXIHP0WCOUNT(),
        .SAXIHP0WDATA(64'd0),
        .SAXIHP0WID(6'd0),
        .SAXIHP0WLAST(1'd0),
        .SAXIHP0WREADY(),
        .SAXIHP0WRISSUECAP1EN(1'd0),
        .SAXIHP0WSTRB(8'd0),
        .SAXIHP0WVALID(1'd0),
        .SAXIHP1ACLK(1'd0),
        .SAXIHP1ARADDR(32'd0),
        .SAXIHP1ARBURST(2'd0),
        .SAXIHP1ARCACHE(4'd0),
        .SAXIHP1ARESETN(),
        .SAXIHP1ARID(6'd0),
        .SAXIHP1ARLEN(4'd0),
        .SAXIHP1ARLOCK(2'd0),
        .SAXIHP1ARPROT(3'd0),
        .SAXIHP1ARQOS(4'd0),
        .SAXIHP1ARREADY(),
        .SAXIHP1ARSIZE(2'd0),
        .SAXIHP1ARVALID(1'd0),
        .SAXIHP1AWADDR(32'd0),
        .SAXIHP1AWBURST(2'd0),
        .SAXIHP1AWCACHE(4'd0),
        .SAXIHP1AWID(6'd0),
        .SAXIHP1AWLEN(4'd0),
        .SAXIHP1AWLOCK(2'd0),
        .SAXIHP1AWPROT(3'd0),
        .SAXIHP1AWQOS(4'd0),
        .SAXIHP1AWREADY(),
        .SAXIHP1AWSIZE(2'd0),
        .SAXIHP1AWVALID(1'd0),
        .SAXIHP1BID(),
        .SAXIHP1BREADY(1'd0),
        .SAXIHP1BRESP(),
        .SAXIHP1BVALID(),
        .SAXIHP1RACOUNT(),
        .SAXIHP1RCOUNT(),
        .SAXIHP1RDATA(),
        .SAXIHP1RDISSUECAP1EN(1'd0),
        .SAXIHP1RID(),
        .SAXIHP1RLAST(),
        .SAXIHP1RREADY(1'd0),
        .SAXIHP1RRESP(),
        .SAXIHP1RVALID(),
        .SAXIHP1WACOUNT(),
        .SAXIHP1WCOUNT(),
        .SAXIHP1WDATA(64'd0),
        .SAXIHP1WID(6'd0),
        .SAXIHP1WLAST(1'd0),
        .SAXIHP1WREADY(),
        .SAXIHP1WRISSUECAP1EN(1'd0),
        .SAXIHP1WSTRB(8'd0),
        .SAXIHP1WVALID(1'd0),
        .SAXIHP2ACLK(1'd0),
        .SAXIHP2ARADDR(32'd0),
        .SAXIHP2ARBURST(2'd0),
        .SAXIHP2ARCACHE(4'd0),
        .SAXIHP2ARESETN(),
        .SAXIHP2ARID(6'd0),
        .SAXIHP2ARLEN(4'd0),
        .SAXIHP2ARLOCK(2'd0),
        .SAXIHP2ARPROT(3'd0),
        .SAXIHP2ARQOS(4'd0),
        .SAXIHP2ARREADY(),
        .SAXIHP2ARSIZE(2'd0),
        .SAXIHP2ARVALID(1'd0),
        .SAXIHP2AWADDR(32'd0),
        .SAXIHP2AWBURST(2'd0),
        .SAXIHP2AWCACHE(4'd0),
        .SAXIHP2AWID(6'd0),
        .SAXIHP2AWLEN(4'd0),
        .SAXIHP2AWLOCK(2'd0),
        .SAXIHP2AWPROT(3'd0),
        .SAXIHP2AWQOS(4'd0),
        .SAXIHP2AWREADY(),
        .SAXIHP2AWSIZE(2'd0),
        .SAXIHP2AWVALID(1'd0),
        .SAXIHP2BID(),
        .SAXIHP2BREADY(1'd0),
        .SAXIHP2BRESP(),
        .SAXIHP2BVALID(),
        .SAXIHP2RACOUNT(),
        .SAXIHP2RCOUNT(),
        .SAXIHP2RDATA(),
        .SAXIHP2RDISSUECAP1EN(1'd0),
        .SAXIHP2RID(),
        .SAXIHP2RLAST(),
        .SAXIHP2RREADY(1'd0),
        .SAXIHP2RRESP(),
        .SAXIHP2RVALID(),
        .SAXIHP2WACOUNT(),
        .SAXIHP2WCOUNT(),
        .SAXIHP2WDATA(64'd0),
        .SAXIHP2WID(6'd0),
        .SAXIHP2WLAST(1'd0),
        .SAXIHP2WREADY(),
        .SAXIHP2WRISSUECAP1EN(1'd0),
        .SAXIHP2WSTRB(8'd0),
        .SAXIHP2WVALID(1'd0),
        .SAXIHP3ACLK(1'd0),
        .SAXIHP3ARADDR(32'd0),
        .SAXIHP3ARBURST(2'd0),
        .SAXIHP3ARCACHE(4'd0),
        .SAXIHP3ARESETN(),
        .SAXIHP3ARID(6'd0),
        .SAXIHP3ARLEN(4'd0),
        .SAXIHP3ARLOCK(2'd0),
        .SAXIHP3ARPROT(3'd0),
        .SAXIHP3ARQOS(4'd0),
        .SAXIHP3ARREADY(),
        .SAXIHP3ARSIZE(2'd0),
        .SAXIHP3ARVALID(1'd0),
        .SAXIHP3AWADDR(32'd0),
        .SAXIHP3AWBURST(2'd0),
        .SAXIHP3AWCACHE(4'd0),
        .SAXIHP3AWID(6'd0),
        .SAXIHP3AWLEN(4'd0),
        .SAXIHP3AWLOCK(2'd0),
        .SAXIHP3AWPROT(3'd0),
        .SAXIHP3AWQOS(4'd0),
        .SAXIHP3AWREADY(),
        .SAXIHP3AWSIZE(2'd0),
        .SAXIHP3AWVALID(1'd0),
        .SAXIHP3BID(),
        .SAXIHP3BREADY(1'd0),
        .SAXIHP3BRESP(),
        .SAXIHP3BVALID(),
        .SAXIHP3RACOUNT(),
        .SAXIHP3RCOUNT(),
        .SAXIHP3RDATA(),
        .SAXIHP3RDISSUECAP1EN(1'd0),
        .SAXIHP3RID(),
        .SAXIHP3RLAST(),
        .SAXIHP3RREADY(1'd0),
        .SAXIHP3RRESP(),
        .SAXIHP3RVALID(),
        .SAXIHP3WACOUNT(),
        .SAXIHP3WCOUNT(),
        .SAXIHP3WDATA(64'd0),
        .SAXIHP3WID(6'd0),
        .SAXIHP3WLAST(1'd0),
        .SAXIHP3WREADY(),
        .SAXIHP3WRISSUECAP1EN(1'd0),
        .SAXIHP3WSTRB(8'd0),
        .SAXIHP3WVALID(1'd0));
    ClockTop pclockTop (
        .CLK(CLK),
        .nRST(nRST),
        .clockOut());
    IOBUF tsda0 (
        .I(pps$EMIOI2C0SDAO),
        .IO(i2c0$sda),
        .O(tsda0$O),
        .T(( !pps$EMIOI2C0SDATN ) && 1'd1));
    IOBUF tscl0 (
        .I(pps$EMIOI2C0SCLO),
        .IO(i2c0$scl),
        .O(tscl0$O),
        .T(( !pps$EMIOI2C0SCLTN ) && 1'd1));
    IOBUF tsda1 (
        .I(pps$EMIOI2C1SDAO),
        .IO(i2c1$sda),
        .O(tsda1$O),
        .T(( !pps$EMIOI2C1SDATN ) && 1'd1));
    IOBUF tscl1 (
        .I(pps$EMIOI2C1SCLO),
        .IO(i2c1$scl),
        .O(tscl1$O),
        .T(( !pps$EMIOI2C1SCLTN ) && 1'd1));
    // Extra assigments, not to output wires
    assign CLK = intr.CLK;
    assign MAXIGP0_O.W$last = pps$MAXIGP0WLAST != 0;
    assign nRST = intr.nRST;
endmodule

`default_nettype wire    // set back to default value
