module PS7 (
  output DMA0DAVALID, output DMA0DRREADY, output DMA0RSTN,
  output DMA1DAVALID, output DMA1DRREADY, output DMA1RSTN,
  output DMA2DAVALID, output DMA2DRREADY, output DMA2RSTN,
  output DMA3DAVALID, output DMA3DRREADY, output DMA3RSTN,
  output EMIOCAN0PHYTX, output EMIOCAN1PHYTX,
  output EMIOENET0GMIITXEN, output EMIOENET0GMIITXER,
  output EMIOENET0MDIOMDC, output EMIOENET0MDIOO, output EMIOENET0MDIOTN,
  output EMIOENET0PTPDELAYREQRX, output EMIOENET0PTPDELAYREQTX,
  output EMIOENET0PTPPDELAYREQRX, output EMIOENET0PTPPDELAYREQTX,
  output EMIOENET0PTPPDELAYRESPRX, output EMIOENET0PTPPDELAYRESPTX,
  output EMIOENET0PTPSYNCFRAMERX, output EMIOENET0PTPSYNCFRAMETX,
  output EMIOENET0SOFRX, output EMIOENET0SOFTX,
  output EMIOENET1GMIITXEN, output EMIOENET1GMIITXER,
  output EMIOENET1MDIOMDC, output EMIOENET1MDIOO, output EMIOENET1MDIOTN,
  output EMIOENET1PTPDELAYREQRX, output EMIOENET1PTPDELAYREQTX,
  output EMIOENET1PTPPDELAYREQRX, output EMIOENET1PTPPDELAYREQTX,
  output EMIOENET1PTPPDELAYRESPRX, output EMIOENET1PTPPDELAYRESPTX,
  output EMIOENET1PTPSYNCFRAMERX, output EMIOENET1PTPSYNCFRAMETX,
  output EMIOENET1SOFRX, output EMIOENET1SOFTX,
  output EMIOI2C0SCLO, output EMIOI2C0SCLTN, output EMIOI2C0SDAO, output EMIOI2C0SDATN,
  output EMIOI2C1SCLO, output EMIOI2C1SCLTN, output EMIOI2C1SDAO, output EMIOI2C1SDATN,
  output EMIOPJTAGTDO, output EMIOPJTAGTDTN,
  output EMIOSDIO0BUSPOW, output EMIOSDIO0CLK, output EMIOSDIO0CMDO, output EMIOSDIO0CMDTN, output EMIOSDIO0LED,
  output EMIOSDIO1BUSPOW, output EMIOSDIO1CLK, output EMIOSDIO1CMDO, output EMIOSDIO1CMDTN, output EMIOSDIO1LED,
  output EMIOSPI0MO, output EMIOSPI0MOTN, output EMIOSPI0SCLKO, output EMIOSPI0SCLKTN,
  output EMIOSPI0SO, output EMIOSPI0SSNTN, output EMIOSPI0STN, output EMIOSPI1MO, output EMIOSPI1MOTN,
  output EMIOSPI1SCLKO, output EMIOSPI1SCLKTN, output EMIOSPI1SO, output EMIOSPI1SSNTN, output EMIOSPI1STN,
  output EMIOTRACECTL,
  output EMIOUART0DTRN, output EMIOUART0RTSN, output EMIOUART0TX,
  output EMIOUART1DTRN, output EMIOUART1RTSN, output EMIOUART1TX,
  output EMIOUSB0VBUSPWRSELECT, output EMIOUSB1VBUSPWRSELECT,
  output EMIOWDTRSTO,
  output EVENTEVENTO,
  output MAXIGP0ARESETN, output MAXIGP0ARVALID, output MAXIGP0AWVALID, output MAXIGP0BREADY, output MAXIGP0RREADY, output MAXIGP0WLAST, output MAXIGP0WVALID,
  output MAXIGP1ARESETN, output MAXIGP1ARVALID, output MAXIGP1AWVALID, output MAXIGP1BREADY, output MAXIGP1RREADY, output MAXIGP1WLAST, output MAXIGP1WVALID,
  output SAXIACPARESETN, output SAXIACPARREADY, output SAXIACPAWREADY, output SAXIACPBVALID, output SAXIACPRLAST, output SAXIACPRVALID, output SAXIACPWREADY,
  output SAXIGP0ARESETN, output SAXIGP0ARREADY, output SAXIGP0AWREADY, output SAXIGP0BVALID, output SAXIGP0RLAST, output SAXIGP0RVALID, output SAXIGP0WREADY,
  output SAXIGP1ARESETN, output SAXIGP1ARREADY, output SAXIGP1AWREADY, output SAXIGP1BVALID, output SAXIGP1RLAST, output SAXIGP1RVALID, output SAXIGP1WREADY,
  output SAXIHP0ARESETN, output SAXIHP0ARREADY, output SAXIHP0AWREADY, output SAXIHP0BVALID, output SAXIHP0RLAST, output SAXIHP0RVALID, output SAXIHP0WREADY,
  output SAXIHP1ARESETN, output SAXIHP1ARREADY, output SAXIHP1AWREADY, output SAXIHP1BVALID, output SAXIHP1RLAST, output SAXIHP1RVALID, output SAXIHP1WREADY,
  output SAXIHP2ARESETN, output SAXIHP2ARREADY, output SAXIHP2AWREADY, output SAXIHP2BVALID, output SAXIHP2RLAST, output SAXIHP2RVALID, output SAXIHP2WREADY,
  output SAXIHP3ARESETN, output SAXIHP3ARREADY, output SAXIHP3AWREADY, output SAXIHP3BVALID, output SAXIHP3RLAST, output SAXIHP3RVALID, output SAXIHP3WREADY,
  output [11:0] MAXIGP0ARID, output [11:0] MAXIGP0AWID, output [11:0] MAXIGP0WID, output [11:0] MAXIGP1ARID, output [11:0] MAXIGP1AWID, output [11:0] MAXIGP1WID,
  output [1:0] DMA0DATYPE, output [1:0] DMA1DATYPE, output [1:0] DMA2DATYPE, output [1:0] DMA3DATYPE,
  output [1:0] EMIOUSB0PORTINDCTL, output [1:0] EMIOUSB1PORTINDCTL,
  output [1:0] EVENTSTANDBYWFE, output [1:0] EVENTSTANDBYWFI,
  output [1:0] MAXIGP0ARBURST, output [1:0] MAXIGP0ARLOCK, output [1:0] MAXIGP0ARSIZE, output [1:0] MAXIGP0AWBURST, output [1:0] MAXIGP0AWLOCK, output [1:0] MAXIGP0AWSIZE,
  output [1:0] MAXIGP1ARBURST, output [1:0] MAXIGP1ARLOCK, output [1:0] MAXIGP1ARSIZE, output [1:0] MAXIGP1AWBURST, output [1:0] MAXIGP1AWLOCK, output [1:0] MAXIGP1AWSIZE,
  output [1:0] SAXIACPBRESP, output [1:0] SAXIACPRRESP,
  output [1:0] SAXIGP0BRESP, output [1:0] SAXIGP0RRESP,
  output [1:0] SAXIGP1BRESP, output [1:0] SAXIGP1RRESP,
  output [1:0] SAXIHP0BRESP, output [1:0] SAXIHP0RRESP,
  output [1:0] SAXIHP1BRESP, output [1:0] SAXIHP1RRESP,
  output [1:0] SAXIHP2BRESP, output [1:0] SAXIHP2RRESP,
  output [1:0] SAXIHP3BRESP, output [1:0] SAXIHP3RRESP,
  output [28:0] IRQP2F,
  output [2:0] EMIOSDIO0BUSVOLT, output [2:0] EMIOSDIO1BUSVOLT,
  output [2:0] EMIOSPI0SSON, output [2:0] EMIOSPI1SSON,
  output [2:0] EMIOTTC0WAVEO, output [2:0] EMIOTTC1WAVEO,
  output [2:0] MAXIGP0ARPROT, output [2:0] MAXIGP0AWPROT,
  output [2:0] MAXIGP1ARPROT, output [2:0] MAXIGP1AWPROT,
  output [2:0] SAXIACPBID, output [2:0] SAXIACPRID,
  output [2:0] SAXIHP0RACOUNT, output [2:0] SAXIHP1RACOUNT, output [2:0] SAXIHP2RACOUNT, output [2:0] SAXIHP3RACOUNT,
  output [31:0] EMIOTRACEDATA,
  output [31:0] FTMTP2FDEBUG,
  output [31:0] MAXIGP0ARADDR, output [31:0] MAXIGP0AWADDR, output [31:0] MAXIGP0WDATA,
  output [31:0] MAXIGP1ARADDR, output [31:0] MAXIGP1AWADDR, output [31:0] MAXIGP1WDATA,
  output [31:0] SAXIGP0RDATA, output [31:0] SAXIGP1RDATA,
  output [3:0] EMIOSDIO0DATAO, output [3:0] EMIOSDIO0DATATN,
  output [3:0] EMIOSDIO1DATAO, output [3:0] EMIOSDIO1DATATN,
  output [3:0] FCLKCLK, output [3:0] FCLKRESETN,
  output [3:0] FTMTF2PTRIGACK, output [3:0] FTMTP2FTRIG,
  output [3:0] MAXIGP0ARCACHE, output [3:0] MAXIGP0ARLEN, output [3:0] MAXIGP0ARQOS, output [3:0] MAXIGP0AWCACHE, output [3:0] MAXIGP0AWLEN, output [3:0] MAXIGP0AWQOS, output [3:0] MAXIGP0WSTRB,
  output [3:0] MAXIGP1ARCACHE, output [3:0] MAXIGP1ARLEN, output [3:0] MAXIGP1ARQOS, output [3:0] MAXIGP1AWCACHE, output [3:0] MAXIGP1AWLEN, output [3:0] MAXIGP1AWQOS, output [3:0] MAXIGP1WSTRB,
  output [5:0] SAXIGP0BID, output [5:0] SAXIGP0RID,
  output [5:0] SAXIGP1BID, output [5:0] SAXIGP1RID,
  output [5:0] SAXIHP0BID, output [5:0] SAXIHP0RID, output [5:0] SAXIHP0WACOUNT,
  output [5:0] SAXIHP1BID, output [5:0] SAXIHP1RID, output [5:0] SAXIHP1WACOUNT,
  output [5:0] SAXIHP2BID, output [5:0] SAXIHP2RID, output [5:0] SAXIHP2WACOUNT,
  output [5:0] SAXIHP3BID, output [5:0] SAXIHP3RID, output [5:0] SAXIHP3WACOUNT,
  output [63:0] EMIOGPIOO, output [63:0] EMIOGPIOTN,
  output [63:0] SAXIACPRDATA, output [63:0] SAXIHP0RDATA, output [63:0] SAXIHP1RDATA, output [63:0] SAXIHP2RDATA, output [63:0] SAXIHP3RDATA,
  output [7:0] EMIOENET0GMIITXD, output [7:0] EMIOENET1GMIITXD,
  output [7:0] SAXIHP0RCOUNT, output [7:0] SAXIHP0WCOUNT,
  output [7:0] SAXIHP1RCOUNT, output [7:0] SAXIHP1WCOUNT,
  output [7:0] SAXIHP2RCOUNT, output [7:0] SAXIHP2WCOUNT,
  output [7:0] SAXIHP3RCOUNT, output [7:0] SAXIHP3WCOUNT,

  inout DDRCASB, inout DDRCKE, inout DDRCKN, inout DDRCKP, inout DDRCSB, inout DDRDRSTB, inout DDRODT, inout DDRRASB, inout DDRVRN, inout DDRVRP, inout DDRWEB,
  inout PSCLK, inout PSPORB, inout PSSRSTB,
  inout [14:0] DDRA, inout [2:0] DDRBA, inout [31:0] DDRDQ, inout [3:0] DDRDM, inout [3:0] DDRDQSN, inout [3:0] DDRDQSP,
  inout [53:0] MIO,
  input DMA0ACLK, input DMA0DAREADY, input DMA0DRLAST, input DMA0DRVALID,
  input DMA1ACLK, input DMA1DAREADY, input DMA1DRLAST, input DMA1DRVALID,
  input DMA2ACLK, input DMA2DAREADY, input DMA2DRLAST, input DMA2DRVALID,
  input DMA3ACLK, input DMA3DAREADY, input DMA3DRLAST, input DMA3DRVALID,
  input EMIOCAN0PHYRX, input EMIOCAN1PHYRX,
  input EMIOENET0EXTINTIN, input EMIOENET0GMIICOL, input EMIOENET0GMIICRS, input EMIOENET0GMIIRXCLK, input EMIOENET0GMIIRXDV, input EMIOENET0GMIIRXER, input EMIOENET0GMIITXCLK, input EMIOENET0MDIOI,
  input EMIOENET1EXTINTIN, input EMIOENET1GMIICOL, input EMIOENET1GMIICRS, input EMIOENET1GMIIRXCLK, input EMIOENET1GMIIRXDV, input EMIOENET1GMIIRXER, input EMIOENET1GMIITXCLK, input EMIOENET1MDIOI,
  input EMIOI2C0SCLI, input EMIOI2C0SDAI,
  input EMIOI2C1SCLI, input EMIOI2C1SDAI,
  input EMIOPJTAGTCK, input EMIOPJTAGTDI, input EMIOPJTAGTMS,
  input EMIOSDIO0CDN, input EMIOSDIO0CLKFB, input EMIOSDIO0CMDI, input EMIOSDIO0WP,
  input EMIOSDIO1CDN, input EMIOSDIO1CLKFB, input EMIOSDIO1CMDI, input EMIOSDIO1WP,
  input EMIOSPI0MI, input EMIOSPI0SCLKI, input EMIOSPI0SI, input EMIOSPI0SSIN,
  input EMIOSPI1MI, input EMIOSPI1SCLKI, input EMIOSPI1SI, input EMIOSPI1SSIN,
  input EMIOSRAMINTIN, input EMIOTRACECLK,
  input EMIOUART0CTSN, input EMIOUART0DCDN, input EMIOUART0DSRN, input EMIOUART0RIN, input EMIOUART0RX,
  input EMIOUART1CTSN, input EMIOUART1DCDN, input EMIOUART1DSRN, input EMIOUART1RIN, input EMIOUART1RX,
  input EMIOUSB0VBUSPWRFAULT, input EMIOUSB1VBUSPWRFAULT,
  input EMIOWDTCLKI,
  input EVENTEVENTI,
  input FPGAIDLEN,
  input FTMDTRACEINCLOCK, input FTMDTRACEINVALID,
  input MAXIGP0ACLK, input MAXIGP0ARREADY, input MAXIGP0AWREADY, input MAXIGP0BVALID, input MAXIGP0RLAST, input MAXIGP0RVALID, input MAXIGP0WREADY,
  input MAXIGP1ACLK, input MAXIGP1ARREADY, input MAXIGP1AWREADY, input MAXIGP1BVALID, input MAXIGP1RLAST, input MAXIGP1RVALID, input MAXIGP1WREADY,
  input SAXIACPACLK, input SAXIACPARVALID, input SAXIACPAWVALID, input SAXIACPBREADY, input SAXIACPRREADY, input SAXIACPWLAST, input SAXIACPWVALID,
  input SAXIGP0ACLK, input SAXIGP0ARVALID, input SAXIGP0AWVALID, input SAXIGP0BREADY, input SAXIGP0RREADY, input SAXIGP0WLAST, input SAXIGP0WVALID,
  input SAXIGP1ACLK, input SAXIGP1ARVALID, input SAXIGP1AWVALID, input SAXIGP1BREADY, input SAXIGP1RREADY, input SAXIGP1WLAST, input SAXIGP1WVALID,
  input SAXIHP0ACLK, input SAXIHP0ARVALID, input SAXIHP0AWVALID, input SAXIHP0BREADY, input SAXIHP0RDISSUECAP1EN, input SAXIHP0RREADY, input SAXIHP0WLAST, input SAXIHP0WRISSUECAP1EN, input SAXIHP0WVALID,
  input SAXIHP1ACLK, input SAXIHP1ARVALID, input SAXIHP1AWVALID, input SAXIHP1BREADY, input SAXIHP1RDISSUECAP1EN, input SAXIHP1RREADY, input SAXIHP1WLAST, input SAXIHP1WRISSUECAP1EN, input SAXIHP1WVALID,
  input SAXIHP2ACLK, input SAXIHP2ARVALID, input SAXIHP2AWVALID, input SAXIHP2BREADY, input SAXIHP2RDISSUECAP1EN, input SAXIHP2RREADY, input SAXIHP2WLAST, input SAXIHP2WRISSUECAP1EN, input SAXIHP2WVALID,
  input SAXIHP3ACLK, input SAXIHP3ARVALID, input SAXIHP3AWVALID, input SAXIHP3BREADY, input SAXIHP3RDISSUECAP1EN, input SAXIHP3RREADY, input SAXIHP3WLAST, input SAXIHP3WRISSUECAP1EN, input SAXIHP3WVALID,
  input [11:0] MAXIGP0BID, input [11:0] MAXIGP0RID,
  input [11:0] MAXIGP1BID, input [11:0] MAXIGP1RID,
  input [19:0] IRQF2P,
  input [1:0] DMA0DRTYPE, input [1:0] DMA1DRTYPE, input [1:0] DMA2DRTYPE, input [1:0] DMA3DRTYPE,
  input [1:0] MAXIGP0BRESP, input [1:0] MAXIGP0RRESP,
  input [1:0] MAXIGP1BRESP, input [1:0] MAXIGP1RRESP,
  input [1:0] SAXIACPARBURST, input [1:0] SAXIACPARLOCK, input [1:0] SAXIACPARSIZE, input [1:0] SAXIACPAWBURST, input [1:0] SAXIACPAWLOCK, input [1:0] SAXIACPAWSIZE,
  input [1:0] SAXIGP0ARBURST, input [1:0] SAXIGP0ARLOCK, input [1:0] SAXIGP0ARSIZE, input [1:0] SAXIGP0AWBURST, input [1:0] SAXIGP0AWLOCK, input [1:0] SAXIGP0AWSIZE,
  input [1:0] SAXIGP1ARBURST, input [1:0] SAXIGP1ARLOCK, input [1:0] SAXIGP1ARSIZE, input [1:0] SAXIGP1AWBURST, input [1:0] SAXIGP1AWLOCK, input [1:0] SAXIGP1AWSIZE,
  input [1:0] SAXIHP0ARBURST, input [1:0] SAXIHP0ARLOCK, input [1:0] SAXIHP0ARSIZE, input [1:0] SAXIHP0AWBURST, input [1:0] SAXIHP0AWLOCK, input [1:0] SAXIHP0AWSIZE,
  input [1:0] SAXIHP1ARBURST, input [1:0] SAXIHP1ARLOCK, input [1:0] SAXIHP1ARSIZE, input [1:0] SAXIHP1AWBURST, input [1:0] SAXIHP1AWLOCK, input [1:0] SAXIHP1AWSIZE,
  input [1:0] SAXIHP2ARBURST, input [1:0] SAXIHP2ARLOCK, input [1:0] SAXIHP2ARSIZE, input [1:0] SAXIHP2AWBURST, input [1:0] SAXIHP2AWLOCK, input [1:0] SAXIHP2AWSIZE,
  input [1:0] SAXIHP3ARBURST, input [1:0] SAXIHP3ARLOCK, input [1:0] SAXIHP3ARSIZE, input [1:0] SAXIHP3AWBURST, input [1:0] SAXIHP3AWLOCK, input [1:0] SAXIHP3AWSIZE,
  input [2:0] EMIOTTC0CLKI, input [2:0] EMIOTTC1CLKI,
  input [2:0] SAXIACPARID, input [2:0] SAXIACPARPROT, input [2:0] SAXIACPAWID, input [2:0] SAXIACPAWPROT, input [2:0] SAXIACPWID,
  input [2:0] SAXIGP0ARPROT, input [2:0] SAXIGP0AWPROT,
  input [2:0] SAXIGP1ARPROT, input [2:0] SAXIGP1AWPROT,
  input [2:0] SAXIHP0ARPROT, input [2:0] SAXIHP0AWPROT,
  input [2:0] SAXIHP1ARPROT, input [2:0] SAXIHP1AWPROT,
  input [2:0] SAXIHP2ARPROT, input [2:0] SAXIHP2AWPROT,
  input [2:0] SAXIHP3ARPROT, input [2:0] SAXIHP3AWPROT,
  input [31:0] FTMDTRACEINDATA, input [31:0] FTMTF2PDEBUG,
  input [31:0] MAXIGP0RDATA, input [31:0] MAXIGP1RDATA,
  input [31:0] SAXIACPARADDR, input [31:0] SAXIACPAWADDR,
  input [31:0] SAXIGP0ARADDR, input [31:0] SAXIGP0AWADDR, input [31:0] SAXIGP0WDATA,
  input [31:0] SAXIGP1ARADDR, input [31:0] SAXIGP1AWADDR, input [31:0] SAXIGP1WDATA,
  input [31:0] SAXIHP0ARADDR, input [31:0] SAXIHP0AWADDR,
  input [31:0] SAXIHP1ARADDR, input [31:0] SAXIHP1AWADDR,
  input [31:0] SAXIHP2ARADDR, input [31:0] SAXIHP2AWADDR,
  input [31:0] SAXIHP3ARADDR, input [31:0] SAXIHP3AWADDR,
  input [3:0] DDRARB,
  input [3:0] EMIOSDIO0DATAI, input [3:0] EMIOSDIO1DATAI,
  input [3:0] FCLKCLKTRIGN,
  input [3:0] FTMDTRACEINATID, input [3:0] FTMTF2PTRIG, input [3:0] FTMTP2FTRIGACK,
  input [3:0] SAXIACPARCACHE, input [3:0] SAXIACPARLEN, input [3:0] SAXIACPARQOS, input [3:0] SAXIACPAWCACHE, input [3:0] SAXIACPAWLEN, input [3:0] SAXIACPAWQOS,
  input [3:0] SAXIGP0ARCACHE, input [3:0] SAXIGP0ARLEN, input [3:0] SAXIGP0ARQOS, input [3:0] SAXIGP0AWCACHE, input [3:0] SAXIGP0AWLEN, input [3:0] SAXIGP0AWQOS, input [3:0] SAXIGP0WSTRB,
  input [3:0] SAXIGP1ARCACHE, input [3:0] SAXIGP1ARLEN, input [3:0] SAXIGP1ARQOS, input [3:0] SAXIGP1AWCACHE, input [3:0] SAXIGP1AWLEN, input [3:0] SAXIGP1AWQOS, input [3:0] SAXIGP1WSTRB,
  input [3:0] SAXIHP0ARCACHE, input [3:0] SAXIHP0ARLEN, input [3:0] SAXIHP0ARQOS, input [3:0] SAXIHP0AWCACHE, input [3:0] SAXIHP0AWLEN, input [3:0] SAXIHP0AWQOS,
  input [3:0] SAXIHP1ARCACHE, input [3:0] SAXIHP1ARLEN, input [3:0] SAXIHP1ARQOS, input [3:0] SAXIHP1AWCACHE, input [3:0] SAXIHP1AWLEN, input [3:0] SAXIHP1AWQOS,
  input [3:0] SAXIHP2ARCACHE, input [3:0] SAXIHP2ARLEN, input [3:0] SAXIHP2ARQOS, input [3:0] SAXIHP2AWCACHE, input [3:0] SAXIHP2AWLEN, input [3:0] SAXIHP2AWQOS,
  input [3:0] SAXIHP3ARCACHE, input [3:0] SAXIHP3ARLEN, input [3:0] SAXIHP3ARQOS, input [3:0] SAXIHP3AWCACHE, input [3:0] SAXIHP3AWLEN, input [3:0] SAXIHP3AWQOS,
  input [4:0] SAXIACPARUSER, input [4:0] SAXIACPAWUSER,
  input [5:0] SAXIGP0ARID, input [5:0] SAXIGP0AWID, input [5:0] SAXIGP0WID,
  input [5:0] SAXIGP1ARID, input [5:0] SAXIGP1AWID, input [5:0] SAXIGP1WID,
  input [5:0] SAXIHP0ARID, input [5:0] SAXIHP0AWID, input [5:0] SAXIHP0WID,
  input [5:0] SAXIHP1ARID, input [5:0] SAXIHP1AWID, input [5:0] SAXIHP1WID,
  input [5:0] SAXIHP2ARID, input [5:0] SAXIHP2AWID, input [5:0] SAXIHP2WID,
  input [5:0] SAXIHP3ARID, input [5:0] SAXIHP3AWID, input [5:0] SAXIHP3WID,
  input [63:0] EMIOGPIOI,
  input [63:0] SAXIACPWDATA, input [63:0] SAXIHP0WDATA, input [63:0] SAXIHP1WDATA, input [63:0] SAXIHP2WDATA, input [63:0] SAXIHP3WDATA,
  input [7:0] EMIOENET0GMIIRXD, input [7:0] EMIOENET1GMIIRXD,
  input [7:0] SAXIACPWSTRB, input [7:0] SAXIHP0WSTRB, input [7:0] SAXIHP1WSTRB, input [7:0] SAXIHP2WSTRB, input [7:0] SAXIHP3WSTRB);
endmodule
