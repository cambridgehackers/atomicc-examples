`ifndef __ft600_GENERATED__VH__
`define __ft600_GENERATED__VH__

//METASTART; ModFt600
//METAINTERNAL; iov; IobufVec;
//METAGUARD; RULE$handshake; 1;
//METARULES; RULE$handshake
`endif
