interface IVectorIndication;
    logic heard__ENA;
    logic [6 - 1:0] heard$meth;
    logic [4 - 1:0] heard$v;
    logic heard__RDY;
    modport server (input  heard__ENA, heard$meth, heard$v,
                    output heard__RDY);
    modport client (output heard__ENA, heard$meth, heard$v,
                    input  heard__RDY);
endinterface
