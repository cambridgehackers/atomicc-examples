`include "atomicclib.vh"

//METASTART; CONNECTNET2
//METAGUARD; RULE$assign; 1'd1;
//METARULES; RULE$assign
