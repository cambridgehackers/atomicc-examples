interface ZynqTopIFC;
    logic [54 - 1:0] MIO;
    logic  I2C0_scl;
    logic  I2C0_sda;
    logic  I2C1_scl;
    logic  I2C1_sda;
endinterface
