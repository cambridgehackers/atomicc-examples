`ifndef __gear1toN_GENERATED__VH__
`define __gear1toN_GENERATED__VH__

//METASTART; Gear1toNBase
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; ( !( 0 == ( ( c == 4 ) ^ 1 ) ) );
//METAGUARD; out$deq; ( !( 0 == ( c == 4 ) ) );
//METAGUARD; out$first; ( !( 0 == ( c == 4 ) ) );
`endif
