`include "atomicclib.vh"

//METASTART; Counter
//METAEXCLUSIVE; startSignal__ENA; RULE$decRule__ENA
//METAGUARD; startSignal; counter == 0;
//METAGUARD; busy; 1'd1;
//METAGUARD; RULE$decRule; counter != 0;
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$decRule; RULE$init
