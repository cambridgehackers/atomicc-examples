
`define BSV_RESET_VALUE 1'b0
`define MAX_IN_WIDTH 128
`define MAX_OUT_WIDTH 128
