`include "atomicclib.vh"

//METASTART; ExternalPin
//METAGUARD; RULE$init; 1'd1;
//METARULES; RULE$init
