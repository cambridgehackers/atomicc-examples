`ifndef __ATOMICCLIB_VH__
`define __ATOMICCLIB_VH__
`include "adapter.generated.vh"
`include "atomicc.generated.vh"
`include "axiTop.generated.vh"
`include "bram.generated.vh"
`include "bscan.generated.vh"
`include "clockTop.generated.vh"
`include "configCounter.generated.vh"
`include "connectNet2.generated.vh"
`include "fifo.generated.vh"
`include "funnel.generated.vh"
`include "grayCounter.generated.vh"
`include "iobufVec.generated.vh"
`include "mimo.generated.vh"
`include "mux.generated.vh"
`include "out2in.generated.vh"
`include "printfStub.generated.vh"
`include "resetInverter.generated.vh"
`include "sizedFifo.generated.vh"
`include "syncFF.generated.vh"
`include "trace.generated.vh"
`include "userTop.generated.vh"
`include "vsimTop.generated.vh"
`include "zynqTop.generated.vh"
`endif
