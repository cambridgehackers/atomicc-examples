`ifndef __asyncControl_GENERATED__VH__
`define __asyncControl_GENERATED__VH__
`include "atomicclib.vh"

//METASTART; AsyncControl
//METAGUARD; RULE$processRule; 1'd1;
//METARULES; RULE$processRule
`endif
