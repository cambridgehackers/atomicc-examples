`ifndef __resetInverter_GENERATED__VH__
`define __resetInverter_GENERATED__VH__

//METASTART; ResetInverter
`endif
