`ifndef __connectNet2_GENERATED__VH__
`define __connectNet2_GENERATED__VH__

//METASTART; CONNECTNET2
//METAGUARD; RULE$assign; 1'd1;
//METARULES; RULE$assign
`endif
