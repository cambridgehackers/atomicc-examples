`include "lpm.generated.vh"

`default_nettype none
module Lpm (input wire CLK, input wire nRST,
    input wire enter__ENA,
    input wire [32 - 1:0]enter$x,
    output wire enter__RDY,
    PipeIn.client outQ);
    ProcessData RULE$enter$agg_2e_tmp;
    wire [32 - 1:0]RULE$enter$x;
    wire RULE$enter__RDY;
    ProcessData RULE$exitr$y;
    wire RULE$exitr__RDY;
    ProcessData RULE$recirc$agg_2e_tmp;
    ProcessData RULE$recirc$y;
    wire RULE$recirc__RDY;
    PipeIn#(.width(23)) fifo$in();
    PipeOut#(.width(23)) fifo$out();
    PipeIn#(.width(32)) inQ$in();
    PipeOut#(.width(32)) inQ$out();
    wire [32 - 1:0]mem$req$v;
    wire mem$req__RDY;
    wire mem$resAccept__RDY;
    wire [32 - 1:0]mem$resValue;
    wire mem$resValue__RDY;
    BufTicket compBuf (.CLK(CLK), .nRST(nRST),
        .getTicket(),
        .getTicket__RDY(),
        .allocateTicket__ENA(0),
        .allocateTicket__RDY());
    Fifo1Base#(.width(32)) inQ (.CLK(CLK), .nRST(nRST),
        .in(inQ$in),
        .out(inQ$out));
    FifoB1Base#(.width(23)) fifo (.CLK(CLK), .nRST(nRST),
        .in(fifo$in),
        .out(fifo$out));
    LpmMemory mem (.CLK(CLK), .nRST(nRST),
        .req__ENA(RULE$recirc__RDY || RULE$enter__RDY),
        .req$v(mem$req$v),
        .req__RDY(mem$req__RDY),
        .resAccept__ENA(RULE$recirc__RDY || RULE$exitr__RDY),
        .resAccept__RDY(mem$resAccept__RDY),
        .resValue(mem$resValue),
        .resValue__RDY(mem$resValue__RDY));
    assign enter__RDY = inQ$in.enq__RDY;
    assign mem$req$v = ( RULE$recirc__RDY ? ( mem$resValue + ( ( RULE$recirc$y.state == 1 ) ? RULE$recirc$y.IPA[ 15 : 8 ] : RULE$recirc$y.IPA[ 7 : 0 ] ) ) : 32'd0 ) | ( RULE$enter__RDY ? ( 32'd0 + RULE$enter$x[ 31 : 16 ] ) : 32'd0 );
    // Extra assigments, not to output wires
    assign RULE$enter$agg_2e_tmp.IPA = RULE$enter$x[ 15 : 0 ];
    assign RULE$enter$agg_2e_tmp.state = 3'd0;
    assign RULE$enter$agg_2e_tmp.ticket = 4'd0;
    assign RULE$enter$x = inQ$out.first;
    assign RULE$enter__RDY = !( ( 0 == ( ( RULE$recirc__RDY != 0 ) ^ 1 ) ) || ( !( inQ$out.first__RDY && inQ$out.deq__RDY && fifo$in.enq__RDY && mem$req__RDY ) ) );
    assign RULE$exitr$y = fifo$out.first;
    assign RULE$exitr__RDY = ( ( mem$resValue & 1 ) == 1 ) && ( RULE$recirc__RDY == 0 ) && mem$resValue__RDY && fifo$out.first__RDY && mem$resAccept__RDY && fifo$out.deq__RDY && outQ.enq__RDY;
    assign RULE$recirc$agg_2e_tmp.IPA = RULE$recirc$y.IPA;
    assign RULE$recirc$agg_2e_tmp.state = RULE$recirc$y.state + 3'd1;
    assign RULE$recirc$agg_2e_tmp.ticket = RULE$recirc$y.ticket;
    assign RULE$recirc$y = fifo$out.first;
    assign RULE$recirc__RDY = !( ( 0 == ( ( ( mem$resValue & 1 ) == 1 ) ^ 1 ) ) || ( !( mem$resValue__RDY && fifo$out.first__RDY && mem$resAccept__RDY && mem$req__RDY && fifo$out.deq__RDY && fifo$in.enq__RDY ) ) );
    assign fifo$in.enq$v = ( RULE$recirc__RDY ? RULE$recirc$agg_2e_tmp : 0 ) | ( RULE$enter__RDY ? RULE$enter$agg_2e_tmp : 0 );
    assign fifo$in.enq__ENA = RULE$recirc__RDY || RULE$enter__RDY;
    assign fifo$out.deq__ENA = RULE$recirc__RDY || RULE$exitr__RDY;
    assign inQ$in.enq$v = enter$x;
    assign inQ$in.enq__ENA = enter__ENA;
    assign inQ$out.deq__ENA = RULE$enter__RDY;
    assign outQ.enq$v = mem$resValue;
    assign outQ.enq__ENA = RULE$exitr__RDY;
endmodule

`default_nettype wire    // set back to default value
