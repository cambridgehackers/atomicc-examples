`ifndef __configCounter_GENERATED__VH__
`define __configCounter_GENERATED__VH__

//METASTART; ConfigCounter
//METAGUARD; RULE$react; 1;
//METAEXCLUSIVE; ifc$decrement__ENA; ifc$maybeDecrement
//METAGUARD; ifc$decrement; 1;
//METAGUARD; ifc$increment; 1;
//METAGUARD; ifc$maybeDecrement; 1;
//METAGUARD; ifc$positive; 1;
//METAGUARD; ifc$read; 1;
//METARULES; RULE$react
`endif
