`ifndef __mimo_GENERATED__VH__
`define __mimo_GENERATED__VH__

//METASTART; MIMOBase
//METAEXCLUSIVE; out$deq__ENA; in$enq__ENA
//METAGUARD; out$deq; c >= widthOut;
//METAGUARD; out$first; c >= widthOut;
//METAGUARD; in$enq; !( c >= widthOut );
`endif
