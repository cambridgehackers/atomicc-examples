`ifndef __configCounter_GENERATED__VH__
`define __configCounter_GENERATED__VH__

//METASTART; ConfigCounter
//METAGUARD; decrement; 1;
//METAGUARD; maybeDecrement; 1;
//METAGUARD; increment; 1;
//METAGUARD; read; 1;
//METAGUARD; positive; 1;
//METAGUARD; RULE$react; 1;
//METARULES; RULE$react
`endif
