`include "hdmi.generated.vh"

`default_nettype none
module HdmiImageon (
    input wire CLK,
    input wire nRST);
endmodule

`default_nettype wire    // set back to default value
