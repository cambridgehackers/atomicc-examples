`ifndef __gear1toN_GENERATED__VH__
`define __gear1toN_GENERATED__VH__

//METASTART; Gear1toNBase
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; c == 0;
//METAGUARD; out$deq; !( c == 0 );
//METAGUARD; out$first; !( c == 0 );
`endif
