`ifndef __funnel_GENERATED__VH__
`define __funnel_GENERATED__VH__

//METASTART; FunnelHalfBase
//METAEXTERNAL; output; FunnelHalfBase$output;
//METAGUARD; input$enq; ( input$enq__ENA[ ( __inst$Genvar1 * 2 ) + 1 ] == 0 ) && output$enq__RDY[ __inst$Genvar1 ];
//METAGUARD; input$enq; input$enq__ENA[ ( __inst$Genvar1 * 2 ) + 1 ] == 0;
`endif
