`ifndef __connectNet2_GENERATED__VH__
`define __connectNet2_GENERATED__VH__

//METASTART; CONNECTNET2
//METAGUARD; RULEassign; 1;
//METARULES; RULEassign
`endif
