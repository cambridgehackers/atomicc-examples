`ifndef __grayCounter_GENERATED__VH__
`define __grayCounter_GENERATED__VH__

//METASTART; GrayCounter
//METAGUARD; RULE$incdec; !( increment__ENA == decrement__ENA );
//METAGUARD; ifc$decrement; 1;
//METAGUARD; ifc$increment; 1;
//METAGUARD; ifc$readBin; 1;
//METAGUARD; ifc$readGray; 1;
//METAGUARD; ifc$writeBin; 1;
//METAGUARD; ifc$writeGray; 1;
//METARULES; RULE$incdec
`endif
