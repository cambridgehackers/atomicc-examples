`ifndef __out2in_GENERATED__VH__
`define __out2in_GENERATED__VH__

//METASTART; Out2In
//METAINVOKE; RULE$copyRule__ENA; :in$deq__ENA;:in$first;:out$enq__ENA;
//METAGUARD; RULE$copyRule; in$first__RDY && out$enq__RDY && in$deq__RDY;
//METARULES; RULE$copyRule
`endif
