`ifndef __iobufVec_GENERATED__VH__
`define __iobufVec_GENERATED__VH__
`include "atomicclib.vh"

`ifndef __IobufVecPins_DEF__
`define __IobufVecPins_DEF__
interface IobufVecPins#(iovecWidth = 999999);
    logic [iovecWidth - 1:0] IO;
    logic [iovecWidth - 1:0] I;
    logic [iovecWidth - 1:0] O;
    logic  T;
    modport server (input  I, T,
                    output O);
    modport client (output I, T,
                    input  O);
endinterface
`endif
//METASTART; IobufVec
//METAINTERNAL; iobufs0; IOBUF;
//METAGUARD; RULE$iobufs; 1;
//METARULES; RULE$iobufs
`endif
