`include "atomicclib.vh"

//METASTART; AsyncControl
//METAGUARD; RULE$processRule; 1'd1;
//METARULES; RULE$processRule
