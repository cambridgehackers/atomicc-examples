`ifndef __before1_GENERATED__VH__
`define __before1_GENERATED__VH__

//METASTART; Connect
//METAEXTERNAL; indication; l_ainterface_OC_EchoIndication;
//METAINTERNAL; lEIO; EchoIndicationOutput;
//METAINTERNAL; lERI; EchoRequestInput;
//METAINTERNAL; lEcho; Echo;
//METAINTERNAL; lERO_test; EchoRequestOutput;
//METAINTERNAL; lEII_test; EchoIndicationInput;
//METAINVOKE; RULEswap2_rule__ENA; :lEcho$swap$y2xnull__ENA;
//METAGUARD; RULEswap2_rule; lEcho$swap$y2xnull__RDY;
//METAINVOKE; RULEswap_rule__ENA; :lEcho$swap$x2y__ENA;:lEcho$swap$y2x__ENA;
//METAGUARD; RULEswap_rule; lEcho$swap$x2y__RDY & lEcho$swap$y2x__RDY;
//METAINVOKE; request$say__ENA; :lERO_test$request$say__ENA;
//METAINVOKE; request$say2__ENA; :lERO_test$request$say2__ENA;
//METAGUARD; request$say2; lERO_test$request$say2__RDY;
//METAGUARD; request$say; lERO_test$request$say__RDY;
//METARULES; RULEswap2_rule; RULEswap_rule
//METACONNECT; lERI$request$say__ENA; lEcho$request$say__ENA
//METACONNECT; lERI$request$say2__ENA; lEcho$request$say2__ENA
//METACONNECT; lERI$request$say2__RDY; lEcho$request$say2__RDY
//METACONNECT; lERI$request$say__RDY; lEcho$request$say__RDY
//METACONNECT; lEIO$pipe$enq__ENA; lEII_test$pipe$enq__ENA
//METACONNECT; lEIO$pipe$enq__RDY; lEII_test$pipe$enq__RDY
//METACONNECT; lEcho$indication$heard__ENA; lEIO$indication$heard__ENA
//METACONNECT; lEcho$indication$heard__RDY; lEIO$indication$heard__RDY
//METACONNECT; lERO_test$pipe$enq__ENA; lERI$pipe$enq__ENA
//METACONNECT; lERO_test$pipe$enq__RDY; lERI$pipe$enq__RDY
//METACONNECT; lEII_test$indication$heard__ENA; indication$heard__ENA
//METACONNECT; lEII_test$indication$heard__RDY; indication$heard__RDY
//METASTART; Echo
//METAEXTERNAL; indication; l_ainterface_OC_EchoIndication;
//METAEXCLUSIVE; RULEdelay_rule__ENA; RULErespond_rule__ENA; request$say2__ENA; request$say__ENA
//METAGUARD; RULEdelay_rule; ( busy & ( !busy_delay ) ) != 0;
//METAINVOKE; RULErespond_rule__ENA; :indication$heard__ENA;
//METAGUARD; RULErespond_rule; busy_delay & indication$heard__RDY;
//METAEXCLUSIVE; request$say__ENA; request$say2__ENA
//METAGUARD; request$say2; !busy;
//METAGUARD; request$say; !busy;
//METAGUARD; swap$x2y; 1;
//METAGUARD; swap$y2x; 1;
//METAGUARD; swap$y2xnull; 1;
//METARULES; RULEdelay_rule; RULErespond_rule
//METASTART; EchoIndicationInput
//METAEXTERNAL; indication; l_ainterface_OC_EchoIndication;
//METAINVOKE; RULEinput_rule__ENA; :indication$heard__ENA;
//METAEXCLUSIVE; RULEinput_rule__ENA; pipe$enq__ENA
//METAGUARD; RULEinput_rule; busy_delay & indication$heard__RDY;
//METAGUARD; pipe$enq; !busy_delay;
//METARULES; RULEinput_rule
//METASTART; EchoIndicationOutput
//METAEXTERNAL; pipe; l_ainterface_OC_PipeIn_OC_1;
//METAINVOKE; RULEoutput_rulee__ENA; :pipe$enq__ENA;
//METAEXCLUSIVE; RULEoutput_rulee__ENA; RULEoutput_ruleo__ENA; indication$heard__ENA
//METAGUARD; RULEoutput_rulee; ( ( ind_busy & even ) != 0 ) & pipe$enq__RDY;
//METAINVOKE; RULEoutput_ruleo__ENA; :pipe$enq__ENA;
//METAEXCLUSIVE; RULEoutput_ruleo__ENA; indication$heard__ENA
//METAGUARD; RULEoutput_ruleo; ( ( ind_busy & ( !even ) ) != 0 ) & pipe$enq__RDY;
//METAGUARD; indication$heard; !ind_busy;
//METARULES; RULEoutput_rulee; RULEoutput_ruleo
//METASTART; EchoRequestInput
//METAEXTERNAL; request; l_ainterface_OC_EchoRequest;
//METAINVOKE; pipe$enq__ENA; pipe$enq__ENA$v_2e_addr$tag == 32'd2:request$say2__ENA;pipe$enq__ENA$v_2e_addr$tag == 32'd1:request$say__ENA;
//METAGUARD; pipe$enq; ( ( pipe$enq__ENA$v_2e_addr$tag != 32'd1 ) | request$say__RDY ) & ( ( pipe$enq__ENA$v_2e_addr$tag != 32'd2 ) | request$say2__RDY );
//METASTART; EchoRequestOutput
//METAEXTERNAL; pipe; l_ainterface_OC_PipeIn_OC_0;
//METAINVOKE; request$say__ENA; :pipe$enq__ENA;
//METAEXCLUSIVE; request$say__ENA; request$say2__ENA
//METAINVOKE; request$say2__ENA; :pipe$enq__ENA;
//METAGUARD; request$say2; pipe$enq__RDY;
//METAGUARD; request$say; pipe$enq__RDY;
//METASTART; Fifo1
//METAEXCLUSIVE; in$enq__ENA; out$deq__ENA
//METAGUARD; in$enq; !full;
//METAGUARD; out$deq; full;
//METAGUARD; out$first; full;
//METASTART; MuxPipe
//METAEXTERNAL; out; l_ainterface_OC_PipeIn;
//METAINTERNAL; forwardFifo; Fifo1;
//METAINVOKE; RULEfifoRule__ENA; :forwardFifo$out$deq__ENA;:forwardFifo$out$first;:out$enq__ENA;
//METAEXCLUSIVE; RULEfifoRule__ENA; in$enq__ENA
//METAGUARD; RULEfifoRule; forwardFifo$out$first__RDY & out$enq__RDY & forwardFifo$out$deq__RDY;
//METAINVOKE; forward$enq__ENA; :forwardFifo$in$enq__ENA;
//METAGUARD; forward$enq; forwardFifo$in$enq__RDY;
//METAINVOKE; in$enq__ENA; :out$enq__ENA;
//METAGUARD; in$enq; out$enq__RDY;
//METARULES; RULEfifoRule
`endif
