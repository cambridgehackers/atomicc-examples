`include "atomicclib.vh"

//METASTART; ModFt600
//METAINTERNAL; iov; IobufVec(iovecWidth=16);
//METAGUARD; RULE$handshake; 1'd1;
//METARULES; RULE$handshake
