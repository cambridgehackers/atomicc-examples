`ifndef __zynqTop_GENERATED__VH__
`define __zynqTop_GENERATED__VH__
`include "atomicclib.vh"

`ifndef __ZynqInterruptT_DEF__
`define __ZynqInterruptT_DEF__
interface ZynqInterruptT;
    logic  CLK;
    logic  nRST;
    logic  interrupt;
    modport server (input  CLK, nRST,
                    output interrupt);
    modport client (output CLK, nRST,
                    input  interrupt);
endinterface
`endif
`ifndef __MaxiO_DEF__
`define __MaxiO_DEF__
interface MaxiO;
    logic AR__ENA;
    logic [32 - 1:0] AR$addr;
    logic [12 - 1:0] AR$id;
    logic [4 - 1:0] AR$len;
    logic AR__RDY;
    logic AW__ENA;
    logic [32 - 1:0] AW$addr;
    logic [12 - 1:0] AW$id;
    logic [4 - 1:0] AW$len;
    logic AW__RDY;
    logic W__ENA;
    logic [32 - 1:0] W$data;
    logic [12 - 1:0] W$id;
    logic  W$last;
    logic W__RDY;
    modport server (input  AR__ENA, AR$addr, AR$id, AR$len, AW__ENA, AW$addr, AW$id, AW$len, W__ENA, W$data, W$id, W$last,
                    output AR__RDY, AW__RDY, W__RDY);
    modport client (output AR__ENA, AR$addr, AR$id, AR$len, AW__ENA, AW$addr, AW$id, AW$len, W__ENA, W$data, W$id, W$last,
                    input  AR__RDY, AW__RDY, W__RDY);
endinterface
`endif
`ifndef __MaxiI_DEF__
`define __MaxiI_DEF__
interface MaxiI;
    logic R__ENA;
    logic [32 - 1:0] R$data;
    logic [12 - 1:0] R$id;
    logic  R$last;
    logic [2 - 1:0] R$resp;
    logic R__RDY;
    logic B__ENA;
    logic [12 - 1:0] B$id;
    logic [2 - 1:0] B$resp;
    logic B__RDY;
    modport server (input  R__ENA, R$data, R$id, R$last, R$resp, B__ENA, B$id, B$resp,
                    output R__RDY, B__RDY);
    modport client (output R__ENA, R$data, R$id, R$last, R$resp, B__ENA, B$id, B$resp,
                    input  R__RDY, B__RDY);
endinterface
`endif
`ifndef __MbufgBUFG_DEF__
`define __MbufgBUFG_DEF__
interface MbufgBUFG;
    logic  I;
    logic  O;
    modport server (input  I,
                    output O);
    modport client (output I,
                    input  O);
endinterface
`endif
`ifndef __ClockIfc_DEF__
`define __ClockIfc_DEF__
interface ClockIfc;
    logic  CLK;
    logic  nRST;
    logic  clockOut;
    modport server (input  CLK, nRST,
                    output clockOut);
    modport client (output CLK, nRST,
                    input  clockOut);
endinterface
`endif
`ifndef __ZynqClock_DEF__
`define __ZynqClock_DEF__
interface ZynqClock;
    logic [15 - 1:0] DDR_Addr;
    logic [3 - 1:0] DDR_BankAddr;
    logic  DDR_CAS_n;
    logic  DDR_CKE;
    logic  DDR_Clk_n;
    logic  DDR_Clk_p;
    logic  DDR_CS_n;
    logic [4 - 1:0] DDR_DM;
    logic [32 - 1:0] DDR_DQ;
    logic [4 - 1:0] DDR_DQS_n;
    logic [4 - 1:0] DDR_DQS_p;
    logic  DDR_DRSTB;
    logic  DDR_ODT;
    logic  DDR_RAS_n;
    logic  FIXED_IO_ddr_vrn;
    logic  FIXED_IO_ddr_vrp;
    logic  DDR_WEB;
    logic  FIXED_IO_ps_clk;
    logic  FIXED_IO_ps_porb;
    logic  FIXED_IO_ps_srstb;
endinterface
`endif
`ifndef __ZynqInterrupt_DEF__
`define __ZynqInterrupt_DEF__
interface ZynqInterrupt;
    logic  interrupt;
    logic  CLK;
    logic  nRST;
    modport server (input  interrupt, CLK, nRST);
    modport client (output interrupt, CLK, nRST);
endinterface
`endif
`ifndef __Pps7fclk_DEF__
`define __Pps7fclk_DEF__
interface Pps7fclk;
    logic [4 - 1:0] CLK;
    logic [4 - 1:0] CLKTRIGN;
    logic [4 - 1:0] RESETN;
    modport server (input  CLKTRIGN,
                    output CLK, RESETN);
    modport client (output CLKTRIGN,
                    input  CLK, RESETN);
endinterface
`endif
`ifndef __P7WrapIfc_DEF__
`define __P7WrapIfc_DEF__
interface P7WrapIfc;
    logic [54 - 1:0] MIO;
endinterface
`endif
`ifndef __Pps7PS7_DEF__
`define __Pps7PS7_DEF__
interface Pps7PS7;
    logic [54 - 1:0] MIO;
    logic [15 - 1:0] DDRA;
    logic [4 - 1:0] DDRARB;
    logic [3 - 1:0] DDRBA;
    logic  DDRCASB;
    logic  DDRCKE;
    logic  DDRCKN;
    logic  DDRCKP;
    logic  DDRCSB;
    logic [4 - 1:0] DDRDM;
    logic [32 - 1:0] DDRDQ;
    logic [4 - 1:0] DDRDQSN;
    logic [4 - 1:0] DDRDQSP;
    logic  DDRDRSTB;
    logic  DDRODT;
    logic  DDRRASB;
    logic  DDRVRN;
    logic  DDRVRP;
    logic  DDRWEB;
    logic  DMA0ACLK;
    logic  DMA0DAREADY;
    logic [2 - 1:0] DMA0DATYPE;
    logic  DMA0DAVALID;
    logic  DMA0DRLAST;
    logic  DMA0DRREADY;
    logic [2 - 1:0] DMA0DRTYPE;
    logic  DMA0DRVALID;
    logic  DMA0RSTN;
    logic  DMA1ACLK;
    logic  DMA1DAREADY;
    logic [2 - 1:0] DMA1DATYPE;
    logic  DMA1DAVALID;
    logic  DMA1DRLAST;
    logic  DMA1DRREADY;
    logic [2 - 1:0] DMA1DRTYPE;
    logic  DMA1DRVALID;
    logic  DMA1RSTN;
    logic  DMA2ACLK;
    logic  DMA2DAREADY;
    logic [2 - 1:0] DMA2DATYPE;
    logic  DMA2DAVALID;
    logic  DMA2DRLAST;
    logic  DMA2DRREADY;
    logic [2 - 1:0] DMA2DRTYPE;
    logic  DMA2DRVALID;
    logic  DMA2RSTN;
    logic  DMA3ACLK;
    logic  DMA3DAREADY;
    logic [2 - 1:0] DMA3DATYPE;
    logic  DMA3DAVALID;
    logic  DMA3DRLAST;
    logic  DMA3DRREADY;
    logic [2 - 1:0] DMA3DRTYPE;
    logic  DMA3DRVALID;
    logic  DMA3RSTN;
    logic  EMIOCAN0PHYRX;
    logic  EMIOCAN0PHYTX;
    logic  EMIOCAN1PHYRX;
    logic  EMIOCAN1PHYTX;
    logic  EMIOENET0EXTINTIN;
    logic  EMIOENET0GMIICOL;
    logic  EMIOENET0GMIICRS;
    logic  EMIOENET0GMIIRXCLK;
    logic [8 - 1:0] EMIOENET0GMIIRXD;
    logic  EMIOENET0GMIIRXDV;
    logic  EMIOENET0GMIIRXER;
    logic  EMIOENET0GMIITXCLK;
    logic [8 - 1:0] EMIOENET0GMIITXD;
    logic  EMIOENET0GMIITXEN;
    logic  EMIOENET0GMIITXER;
    logic  EMIOENET0MDIOI;
    logic  EMIOENET0MDIOMDC;
    logic  EMIOENET0MDIOO;
    logic  EMIOENET0MDIOTN;
    logic  EMIOENET0PTPDELAYREQRX;
    logic  EMIOENET0PTPDELAYREQTX;
    logic  EMIOENET0PTPPDELAYREQRX;
    logic  EMIOENET0PTPPDELAYREQTX;
    logic  EMIOENET0PTPPDELAYRESPRX;
    logic  EMIOENET0PTPPDELAYRESPTX;
    logic  EMIOENET0PTPSYNCFRAMERX;
    logic  EMIOENET0PTPSYNCFRAMETX;
    logic  EMIOENET0SOFRX;
    logic  EMIOENET0SOFTX;
    logic  EMIOENET1EXTINTIN;
    logic  EMIOENET1GMIICOL;
    logic  EMIOENET1GMIICRS;
    logic  EMIOENET1GMIIRXCLK;
    logic [8 - 1:0] EMIOENET1GMIIRXD;
    logic  EMIOENET1GMIIRXDV;
    logic  EMIOENET1GMIIRXER;
    logic  EMIOENET1GMIITXCLK;
    logic [8 - 1:0] EMIOENET1GMIITXD;
    logic  EMIOENET1GMIITXEN;
    logic  EMIOENET1GMIITXER;
    logic  EMIOENET1MDIOI;
    logic  EMIOENET1MDIOMDC;
    logic  EMIOENET1MDIOO;
    logic  EMIOENET1MDIOTN;
    logic  EMIOENET1PTPDELAYREQRX;
    logic  EMIOENET1PTPDELAYREQTX;
    logic  EMIOENET1PTPPDELAYREQRX;
    logic  EMIOENET1PTPPDELAYREQTX;
    logic  EMIOENET1PTPPDELAYRESPRX;
    logic  EMIOENET1PTPPDELAYRESPTX;
    logic  EMIOENET1PTPSYNCFRAMERX;
    logic  EMIOENET1PTPSYNCFRAMETX;
    logic  EMIOENET1SOFRX;
    logic  EMIOENET1SOFTX;
    logic [64 - 1:0] EMIOGPIOI;
    logic [64 - 1:0] EMIOGPIOO;
    logic [64 - 1:0] EMIOGPIOTN;
    logic  EMIOI2C0SCLI;
    logic  EMIOI2C0SCLO;
    logic  EMIOI2C0SCLTN;
    logic  EMIOI2C0SDAI;
    logic  EMIOI2C0SDAO;
    logic  EMIOI2C0SDATN;
    logic  EMIOI2C1SCLI;
    logic  EMIOI2C1SCLO;
    logic  EMIOI2C1SCLTN;
    logic  EMIOI2C1SDAI;
    logic  EMIOI2C1SDAO;
    logic  EMIOI2C1SDATN;
    logic  EMIOPJTAGTCK;
    logic  EMIOPJTAGTDI;
    logic  EMIOPJTAGTDO;
    logic  EMIOPJTAGTDTN;
    logic  EMIOPJTAGTMS;
    logic  EMIOSDIO0BUSPOW;
    logic [3 - 1:0] EMIOSDIO0BUSVOLT;
    logic  EMIOSDIO0CDN;
    logic  EMIOSDIO0CLK;
    logic  EMIOSDIO0CLKFB;
    logic  EMIOSDIO0CMDI;
    logic  EMIOSDIO0CMDO;
    logic  EMIOSDIO0CMDTN;
    logic [4 - 1:0] EMIOSDIO0DATAI;
    logic [4 - 1:0] EMIOSDIO0DATAO;
    logic [4 - 1:0] EMIOSDIO0DATATN;
    logic  EMIOSDIO0LED;
    logic  EMIOSDIO0WP;
    logic  EMIOSDIO1BUSPOW;
    logic [3 - 1:0] EMIOSDIO1BUSVOLT;
    logic  EMIOSDIO1CDN;
    logic  EMIOSDIO1CLK;
    logic  EMIOSDIO1CLKFB;
    logic  EMIOSDIO1CMDI;
    logic  EMIOSDIO1CMDO;
    logic  EMIOSDIO1CMDTN;
    logic [4 - 1:0] EMIOSDIO1DATAI;
    logic [4 - 1:0] EMIOSDIO1DATAO;
    logic [4 - 1:0] EMIOSDIO1DATATN;
    logic  EMIOSDIO1LED;
    logic  EMIOSDIO1WP;
    logic  EMIOSPI0MI;
    logic  EMIOSPI0MO;
    logic  EMIOSPI0MOTN;
    logic  EMIOSPI0SCLKI;
    logic  EMIOSPI0SCLKO;
    logic  EMIOSPI0SCLKTN;
    logic  EMIOSPI0SI;
    logic  EMIOSPI0SO;
    logic  EMIOSPI0SSIN;
    logic  EMIOSPI0SSNTN;
    logic [3 - 1:0] EMIOSPI0SSON;
    logic  EMIOSPI0STN;
    logic  EMIOSPI1MI;
    logic  EMIOSPI1MO;
    logic  EMIOSPI1MOTN;
    logic  EMIOSPI1SCLKI;
    logic  EMIOSPI1SCLKO;
    logic  EMIOSPI1SCLKTN;
    logic  EMIOSPI1SI;
    logic  EMIOSPI1SO;
    logic  EMIOSPI1SSIN;
    logic  EMIOSPI1SSNTN;
    logic [3 - 1:0] EMIOSPI1SSON;
    logic  EMIOSPI1STN;
    logic  EMIOSRAMINTIN;
    logic  EMIOTRACECLK;
    logic  EMIOTRACECTL;
    logic [32 - 1:0] EMIOTRACEDATA;
    logic [3 - 1:0] EMIOTTC0CLKI;
    logic [3 - 1:0] EMIOTTC0WAVEO;
    logic [3 - 1:0] EMIOTTC1CLKI;
    logic [3 - 1:0] EMIOTTC1WAVEO;
    logic  EMIOUART0CTSN;
    logic  EMIOUART0DCDN;
    logic  EMIOUART0DSRN;
    logic  EMIOUART0DTRN;
    logic  EMIOUART0RIN;
    logic  EMIOUART0RTSN;
    logic  EMIOUART0RX;
    logic  EMIOUART0TX;
    logic  EMIOUART1CTSN;
    logic  EMIOUART1DCDN;
    logic  EMIOUART1DSRN;
    logic  EMIOUART1DTRN;
    logic  EMIOUART1RIN;
    logic  EMIOUART1RTSN;
    logic  EMIOUART1RX;
    logic  EMIOUART1TX;
    logic [2 - 1:0] EMIOUSB0PORTINDCTL;
    logic  EMIOUSB0VBUSPWRFAULT;
    logic  EMIOUSB0VBUSPWRSELECT;
    logic [2 - 1:0] EMIOUSB1PORTINDCTL;
    logic  EMIOUSB1VBUSPWRFAULT;
    logic  EMIOUSB1VBUSPWRSELECT;
    logic  EMIOWDTCLKI;
    logic  EMIOWDTRSTO;
    logic  EVENTEVENTI;
    logic  EVENTEVENTO;
    logic [2 - 1:0] EVENTSTANDBYWFE;
    logic [2 - 1:0] EVENTSTANDBYWFI;
    logic [4 - 1:0] FCLKCLK;
    logic [4 - 1:0] FCLKCLKTRIGN;
    logic [4 - 1:0] FCLKRESETN;
    logic  FPGAIDLEN;
    logic [4 - 1:0] FTMDTRACEINATID;
    logic  FTMDTRACEINCLOCK;
    logic [32 - 1:0] FTMDTRACEINDATA;
    logic  FTMDTRACEINVALID;
    logic [32 - 1:0] FTMTF2PDEBUG;
    logic [4 - 1:0] FTMTF2PTRIG;
    logic [4 - 1:0] FTMTF2PTRIGACK;
    logic [32 - 1:0] FTMTP2FDEBUG;
    logic [4 - 1:0] FTMTP2FTRIG;
    logic [4 - 1:0] FTMTP2FTRIGACK;
    logic [20 - 1:0] IRQF2P;
    logic [29 - 1:0] IRQP2F;
    logic  MAXIGP0ACLK;
    logic [32 - 1:0] MAXIGP0ARADDR;
    logic [2 - 1:0] MAXIGP0ARBURST;
    logic [4 - 1:0] MAXIGP0ARCACHE;
    logic  MAXIGP0ARESETN;
    logic [12 - 1:0] MAXIGP0ARID;
    logic [4 - 1:0] MAXIGP0ARLEN;
    logic [2 - 1:0] MAXIGP0ARLOCK;
    logic [3 - 1:0] MAXIGP0ARPROT;
    logic [4 - 1:0] MAXIGP0ARQOS;
    logic  MAXIGP0ARREADY;
    logic [2 - 1:0] MAXIGP0ARSIZE;
    logic  MAXIGP0ARVALID;
    logic [32 - 1:0] MAXIGP0AWADDR;
    logic [2 - 1:0] MAXIGP0AWBURST;
    logic [4 - 1:0] MAXIGP0AWCACHE;
    logic [12 - 1:0] MAXIGP0AWID;
    logic [4 - 1:0] MAXIGP0AWLEN;
    logic [2 - 1:0] MAXIGP0AWLOCK;
    logic [3 - 1:0] MAXIGP0AWPROT;
    logic [4 - 1:0] MAXIGP0AWQOS;
    logic  MAXIGP0AWREADY;
    logic [2 - 1:0] MAXIGP0AWSIZE;
    logic  MAXIGP0AWVALID;
    logic [12 - 1:0] MAXIGP0BID;
    logic  MAXIGP0BREADY;
    logic [2 - 1:0] MAXIGP0BRESP;
    logic  MAXIGP0BVALID;
    logic [32 - 1:0] MAXIGP0RDATA;
    logic [12 - 1:0] MAXIGP0RID;
    logic  MAXIGP0RLAST;
    logic  MAXIGP0RREADY;
    logic [2 - 1:0] MAXIGP0RRESP;
    logic  MAXIGP0RVALID;
    logic [32 - 1:0] MAXIGP0WDATA;
    logic [12 - 1:0] MAXIGP0WID;
    logic  MAXIGP0WLAST;
    logic  MAXIGP0WREADY;
    logic [4 - 1:0] MAXIGP0WSTRB;
    logic  MAXIGP0WVALID;
    logic  MAXIGP1ACLK;
    logic [32 - 1:0] MAXIGP1ARADDR;
    logic [2 - 1:0] MAXIGP1ARBURST;
    logic [4 - 1:0] MAXIGP1ARCACHE;
    logic  MAXIGP1ARESETN;
    logic [12 - 1:0] MAXIGP1ARID;
    logic [4 - 1:0] MAXIGP1ARLEN;
    logic [2 - 1:0] MAXIGP1ARLOCK;
    logic [3 - 1:0] MAXIGP1ARPROT;
    logic [4 - 1:0] MAXIGP1ARQOS;
    logic  MAXIGP1ARREADY;
    logic [2 - 1:0] MAXIGP1ARSIZE;
    logic  MAXIGP1ARVALID;
    logic [32 - 1:0] MAXIGP1AWADDR;
    logic [2 - 1:0] MAXIGP1AWBURST;
    logic [4 - 1:0] MAXIGP1AWCACHE;
    logic [12 - 1:0] MAXIGP1AWID;
    logic [4 - 1:0] MAXIGP1AWLEN;
    logic [2 - 1:0] MAXIGP1AWLOCK;
    logic [3 - 1:0] MAXIGP1AWPROT;
    logic [4 - 1:0] MAXIGP1AWQOS;
    logic  MAXIGP1AWREADY;
    logic [2 - 1:0] MAXIGP1AWSIZE;
    logic  MAXIGP1AWVALID;
    logic [12 - 1:0] MAXIGP1BID;
    logic  MAXIGP1BREADY;
    logic [2 - 1:0] MAXIGP1BRESP;
    logic  MAXIGP1BVALID;
    logic [32 - 1:0] MAXIGP1RDATA;
    logic [12 - 1:0] MAXIGP1RID;
    logic  MAXIGP1RLAST;
    logic  MAXIGP1RREADY;
    logic [2 - 1:0] MAXIGP1RRESP;
    logic  MAXIGP1RVALID;
    logic [32 - 1:0] MAXIGP1WDATA;
    logic [12 - 1:0] MAXIGP1WID;
    logic  MAXIGP1WLAST;
    logic  MAXIGP1WREADY;
    logic [4 - 1:0] MAXIGP1WSTRB;
    logic  MAXIGP1WVALID;
    logic  PSCLK;
    logic  PSPORB;
    logic  PSSRSTB;
    logic  SAXIACPACLK;
    logic [32 - 1:0] SAXIACPARADDR;
    logic [2 - 1:0] SAXIACPARBURST;
    logic [4 - 1:0] SAXIACPARCACHE;
    logic  SAXIACPARESETN;
    logic [3 - 1:0] SAXIACPARID;
    logic [4 - 1:0] SAXIACPARLEN;
    logic [2 - 1:0] SAXIACPARLOCK;
    logic [3 - 1:0] SAXIACPARPROT;
    logic [4 - 1:0] SAXIACPARQOS;
    logic  SAXIACPARREADY;
    logic [2 - 1:0] SAXIACPARSIZE;
    logic [5 - 1:0] SAXIACPARUSER;
    logic  SAXIACPARVALID;
    logic [32 - 1:0] SAXIACPAWADDR;
    logic [2 - 1:0] SAXIACPAWBURST;
    logic [4 - 1:0] SAXIACPAWCACHE;
    logic [3 - 1:0] SAXIACPAWID;
    logic [4 - 1:0] SAXIACPAWLEN;
    logic [2 - 1:0] SAXIACPAWLOCK;
    logic [3 - 1:0] SAXIACPAWPROT;
    logic [4 - 1:0] SAXIACPAWQOS;
    logic  SAXIACPAWREADY;
    logic [2 - 1:0] SAXIACPAWSIZE;
    logic [5 - 1:0] SAXIACPAWUSER;
    logic  SAXIACPAWVALID;
    logic [3 - 1:0] SAXIACPBID;
    logic  SAXIACPBREADY;
    logic [2 - 1:0] SAXIACPBRESP;
    logic  SAXIACPBVALID;
    logic [64 - 1:0] SAXIACPRDATA;
    logic [3 - 1:0] SAXIACPRID;
    logic  SAXIACPRLAST;
    logic  SAXIACPRREADY;
    logic [2 - 1:0] SAXIACPRRESP;
    logic  SAXIACPRVALID;
    logic [64 - 1:0] SAXIACPWDATA;
    logic [3 - 1:0] SAXIACPWID;
    logic  SAXIACPWLAST;
    logic  SAXIACPWREADY;
    logic [8 - 1:0] SAXIACPWSTRB;
    logic  SAXIACPWVALID;
    logic  SAXIGP0ACLK;
    logic [32 - 1:0] SAXIGP0ARADDR;
    logic [2 - 1:0] SAXIGP0ARBURST;
    logic [4 - 1:0] SAXIGP0ARCACHE;
    logic  SAXIGP0ARESETN;
    logic [6 - 1:0] SAXIGP0ARID;
    logic [4 - 1:0] SAXIGP0ARLEN;
    logic [2 - 1:0] SAXIGP0ARLOCK;
    logic [3 - 1:0] SAXIGP0ARPROT;
    logic [4 - 1:0] SAXIGP0ARQOS;
    logic  SAXIGP0ARREADY;
    logic [2 - 1:0] SAXIGP0ARSIZE;
    logic  SAXIGP0ARVALID;
    logic [32 - 1:0] SAXIGP0AWADDR;
    logic [2 - 1:0] SAXIGP0AWBURST;
    logic [4 - 1:0] SAXIGP0AWCACHE;
    logic [6 - 1:0] SAXIGP0AWID;
    logic [4 - 1:0] SAXIGP0AWLEN;
    logic [2 - 1:0] SAXIGP0AWLOCK;
    logic [3 - 1:0] SAXIGP0AWPROT;
    logic [4 - 1:0] SAXIGP0AWQOS;
    logic  SAXIGP0AWREADY;
    logic [2 - 1:0] SAXIGP0AWSIZE;
    logic  SAXIGP0AWVALID;
    logic [6 - 1:0] SAXIGP0BID;
    logic  SAXIGP0BREADY;
    logic [2 - 1:0] SAXIGP0BRESP;
    logic  SAXIGP0BVALID;
    logic [32 - 1:0] SAXIGP0RDATA;
    logic [6 - 1:0] SAXIGP0RID;
    logic  SAXIGP0RLAST;
    logic  SAXIGP0RREADY;
    logic [2 - 1:0] SAXIGP0RRESP;
    logic  SAXIGP0RVALID;
    logic [32 - 1:0] SAXIGP0WDATA;
    logic [6 - 1:0] SAXIGP0WID;
    logic  SAXIGP0WLAST;
    logic  SAXIGP0WREADY;
    logic [4 - 1:0] SAXIGP0WSTRB;
    logic  SAXIGP0WVALID;
    logic  SAXIGP1ACLK;
    logic [32 - 1:0] SAXIGP1ARADDR;
    logic [2 - 1:0] SAXIGP1ARBURST;
    logic [4 - 1:0] SAXIGP1ARCACHE;
    logic  SAXIGP1ARESETN;
    logic [6 - 1:0] SAXIGP1ARID;
    logic [4 - 1:0] SAXIGP1ARLEN;
    logic [2 - 1:0] SAXIGP1ARLOCK;
    logic [3 - 1:0] SAXIGP1ARPROT;
    logic [4 - 1:0] SAXIGP1ARQOS;
    logic  SAXIGP1ARREADY;
    logic [2 - 1:0] SAXIGP1ARSIZE;
    logic  SAXIGP1ARVALID;
    logic [32 - 1:0] SAXIGP1AWADDR;
    logic [2 - 1:0] SAXIGP1AWBURST;
    logic [4 - 1:0] SAXIGP1AWCACHE;
    logic [6 - 1:0] SAXIGP1AWID;
    logic [4 - 1:0] SAXIGP1AWLEN;
    logic [2 - 1:0] SAXIGP1AWLOCK;
    logic [3 - 1:0] SAXIGP1AWPROT;
    logic [4 - 1:0] SAXIGP1AWQOS;
    logic  SAXIGP1AWREADY;
    logic [2 - 1:0] SAXIGP1AWSIZE;
    logic  SAXIGP1AWVALID;
    logic [6 - 1:0] SAXIGP1BID;
    logic  SAXIGP1BREADY;
    logic [2 - 1:0] SAXIGP1BRESP;
    logic  SAXIGP1BVALID;
    logic [32 - 1:0] SAXIGP1RDATA;
    logic [6 - 1:0] SAXIGP1RID;
    logic  SAXIGP1RLAST;
    logic  SAXIGP1RREADY;
    logic [2 - 1:0] SAXIGP1RRESP;
    logic  SAXIGP1RVALID;
    logic [32 - 1:0] SAXIGP1WDATA;
    logic [6 - 1:0] SAXIGP1WID;
    logic  SAXIGP1WLAST;
    logic  SAXIGP1WREADY;
    logic [4 - 1:0] SAXIGP1WSTRB;
    logic  SAXIGP1WVALID;
    logic  SAXIHP0ACLK;
    logic [32 - 1:0] SAXIHP0ARADDR;
    logic [2 - 1:0] SAXIHP0ARBURST;
    logic [4 - 1:0] SAXIHP0ARCACHE;
    logic  SAXIHP0ARESETN;
    logic [6 - 1:0] SAXIHP0ARID;
    logic [4 - 1:0] SAXIHP0ARLEN;
    logic [2 - 1:0] SAXIHP0ARLOCK;
    logic [3 - 1:0] SAXIHP0ARPROT;
    logic [4 - 1:0] SAXIHP0ARQOS;
    logic  SAXIHP0ARREADY;
    logic [2 - 1:0] SAXIHP0ARSIZE;
    logic  SAXIHP0ARVALID;
    logic [32 - 1:0] SAXIHP0AWADDR;
    logic [2 - 1:0] SAXIHP0AWBURST;
    logic [4 - 1:0] SAXIHP0AWCACHE;
    logic [6 - 1:0] SAXIHP0AWID;
    logic [4 - 1:0] SAXIHP0AWLEN;
    logic [2 - 1:0] SAXIHP0AWLOCK;
    logic [3 - 1:0] SAXIHP0AWPROT;
    logic [4 - 1:0] SAXIHP0AWQOS;
    logic  SAXIHP0AWREADY;
    logic [2 - 1:0] SAXIHP0AWSIZE;
    logic  SAXIHP0AWVALID;
    logic [6 - 1:0] SAXIHP0BID;
    logic  SAXIHP0BREADY;
    logic [2 - 1:0] SAXIHP0BRESP;
    logic  SAXIHP0BVALID;
    logic [3 - 1:0] SAXIHP0RACOUNT;
    logic [8 - 1:0] SAXIHP0RCOUNT;
    logic [64 - 1:0] SAXIHP0RDATA;
    logic  SAXIHP0RDISSUECAP1EN;
    logic [6 - 1:0] SAXIHP0RID;
    logic  SAXIHP0RLAST;
    logic  SAXIHP0RREADY;
    logic [2 - 1:0] SAXIHP0RRESP;
    logic  SAXIHP0RVALID;
    logic [6 - 1:0] SAXIHP0WACOUNT;
    logic [8 - 1:0] SAXIHP0WCOUNT;
    logic [64 - 1:0] SAXIHP0WDATA;
    logic [6 - 1:0] SAXIHP0WID;
    logic  SAXIHP0WLAST;
    logic  SAXIHP0WREADY;
    logic  SAXIHP0WRISSUECAP1EN;
    logic [8 - 1:0] SAXIHP0WSTRB;
    logic  SAXIHP0WVALID;
    logic  SAXIHP1ACLK;
    logic [32 - 1:0] SAXIHP1ARADDR;
    logic [2 - 1:0] SAXIHP1ARBURST;
    logic [4 - 1:0] SAXIHP1ARCACHE;
    logic  SAXIHP1ARESETN;
    logic [6 - 1:0] SAXIHP1ARID;
    logic [4 - 1:0] SAXIHP1ARLEN;
    logic [2 - 1:0] SAXIHP1ARLOCK;
    logic [3 - 1:0] SAXIHP1ARPROT;
    logic [4 - 1:0] SAXIHP1ARQOS;
    logic  SAXIHP1ARREADY;
    logic [2 - 1:0] SAXIHP1ARSIZE;
    logic  SAXIHP1ARVALID;
    logic [32 - 1:0] SAXIHP1AWADDR;
    logic [2 - 1:0] SAXIHP1AWBURST;
    logic [4 - 1:0] SAXIHP1AWCACHE;
    logic [6 - 1:0] SAXIHP1AWID;
    logic [4 - 1:0] SAXIHP1AWLEN;
    logic [2 - 1:0] SAXIHP1AWLOCK;
    logic [3 - 1:0] SAXIHP1AWPROT;
    logic [4 - 1:0] SAXIHP1AWQOS;
    logic  SAXIHP1AWREADY;
    logic [2 - 1:0] SAXIHP1AWSIZE;
    logic  SAXIHP1AWVALID;
    logic [6 - 1:0] SAXIHP1BID;
    logic  SAXIHP1BREADY;
    logic [2 - 1:0] SAXIHP1BRESP;
    logic  SAXIHP1BVALID;
    logic [3 - 1:0] SAXIHP1RACOUNT;
    logic [8 - 1:0] SAXIHP1RCOUNT;
    logic [64 - 1:0] SAXIHP1RDATA;
    logic  SAXIHP1RDISSUECAP1EN;
    logic [6 - 1:0] SAXIHP1RID;
    logic  SAXIHP1RLAST;
    logic  SAXIHP1RREADY;
    logic [2 - 1:0] SAXIHP1RRESP;
    logic  SAXIHP1RVALID;
    logic [6 - 1:0] SAXIHP1WACOUNT;
    logic [8 - 1:0] SAXIHP1WCOUNT;
    logic [64 - 1:0] SAXIHP1WDATA;
    logic [6 - 1:0] SAXIHP1WID;
    logic  SAXIHP1WLAST;
    logic  SAXIHP1WREADY;
    logic  SAXIHP1WRISSUECAP1EN;
    logic [8 - 1:0] SAXIHP1WSTRB;
    logic  SAXIHP1WVALID;
    logic  SAXIHP2ACLK;
    logic [32 - 1:0] SAXIHP2ARADDR;
    logic [2 - 1:0] SAXIHP2ARBURST;
    logic [4 - 1:0] SAXIHP2ARCACHE;
    logic  SAXIHP2ARESETN;
    logic [6 - 1:0] SAXIHP2ARID;
    logic [4 - 1:0] SAXIHP2ARLEN;
    logic [2 - 1:0] SAXIHP2ARLOCK;
    logic [3 - 1:0] SAXIHP2ARPROT;
    logic [4 - 1:0] SAXIHP2ARQOS;
    logic  SAXIHP2ARREADY;
    logic [2 - 1:0] SAXIHP2ARSIZE;
    logic  SAXIHP2ARVALID;
    logic [32 - 1:0] SAXIHP2AWADDR;
    logic [2 - 1:0] SAXIHP2AWBURST;
    logic [4 - 1:0] SAXIHP2AWCACHE;
    logic [6 - 1:0] SAXIHP2AWID;
    logic [4 - 1:0] SAXIHP2AWLEN;
    logic [2 - 1:0] SAXIHP2AWLOCK;
    logic [3 - 1:0] SAXIHP2AWPROT;
    logic [4 - 1:0] SAXIHP2AWQOS;
    logic  SAXIHP2AWREADY;
    logic [2 - 1:0] SAXIHP2AWSIZE;
    logic  SAXIHP2AWVALID;
    logic [6 - 1:0] SAXIHP2BID;
    logic  SAXIHP2BREADY;
    logic [2 - 1:0] SAXIHP2BRESP;
    logic  SAXIHP2BVALID;
    logic [3 - 1:0] SAXIHP2RACOUNT;
    logic [8 - 1:0] SAXIHP2RCOUNT;
    logic [64 - 1:0] SAXIHP2RDATA;
    logic  SAXIHP2RDISSUECAP1EN;
    logic [6 - 1:0] SAXIHP2RID;
    logic  SAXIHP2RLAST;
    logic  SAXIHP2RREADY;
    logic [2 - 1:0] SAXIHP2RRESP;
    logic  SAXIHP2RVALID;
    logic [6 - 1:0] SAXIHP2WACOUNT;
    logic [8 - 1:0] SAXIHP2WCOUNT;
    logic [64 - 1:0] SAXIHP2WDATA;
    logic [6 - 1:0] SAXIHP2WID;
    logic  SAXIHP2WLAST;
    logic  SAXIHP2WREADY;
    logic  SAXIHP2WRISSUECAP1EN;
    logic [8 - 1:0] SAXIHP2WSTRB;
    logic  SAXIHP2WVALID;
    logic  SAXIHP3ACLK;
    logic [32 - 1:0] SAXIHP3ARADDR;
    logic [2 - 1:0] SAXIHP3ARBURST;
    logic [4 - 1:0] SAXIHP3ARCACHE;
    logic  SAXIHP3ARESETN;
    logic [6 - 1:0] SAXIHP3ARID;
    logic [4 - 1:0] SAXIHP3ARLEN;
    logic [2 - 1:0] SAXIHP3ARLOCK;
    logic [3 - 1:0] SAXIHP3ARPROT;
    logic [4 - 1:0] SAXIHP3ARQOS;
    logic  SAXIHP3ARREADY;
    logic [2 - 1:0] SAXIHP3ARSIZE;
    logic  SAXIHP3ARVALID;
    logic [32 - 1:0] SAXIHP3AWADDR;
    logic [2 - 1:0] SAXIHP3AWBURST;
    logic [4 - 1:0] SAXIHP3AWCACHE;
    logic [6 - 1:0] SAXIHP3AWID;
    logic [4 - 1:0] SAXIHP3AWLEN;
    logic [2 - 1:0] SAXIHP3AWLOCK;
    logic [3 - 1:0] SAXIHP3AWPROT;
    logic [4 - 1:0] SAXIHP3AWQOS;
    logic  SAXIHP3AWREADY;
    logic [2 - 1:0] SAXIHP3AWSIZE;
    logic  SAXIHP3AWVALID;
    logic [6 - 1:0] SAXIHP3BID;
    logic  SAXIHP3BREADY;
    logic [2 - 1:0] SAXIHP3BRESP;
    logic  SAXIHP3BVALID;
    logic [3 - 1:0] SAXIHP3RACOUNT;
    logic [8 - 1:0] SAXIHP3RCOUNT;
    logic [64 - 1:0] SAXIHP3RDATA;
    logic  SAXIHP3RDISSUECAP1EN;
    logic [6 - 1:0] SAXIHP3RID;
    logic  SAXIHP3RLAST;
    logic  SAXIHP3RREADY;
    logic [2 - 1:0] SAXIHP3RRESP;
    logic  SAXIHP3RVALID;
    logic [6 - 1:0] SAXIHP3WACOUNT;
    logic [8 - 1:0] SAXIHP3WCOUNT;
    logic [64 - 1:0] SAXIHP3WDATA;
    logic [6 - 1:0] SAXIHP3WID;
    logic  SAXIHP3WLAST;
    logic  SAXIHP3WREADY;
    logic  SAXIHP3WRISSUECAP1EN;
    logic [8 - 1:0] SAXIHP3WSTRB;
    logic  SAXIHP3WVALID;
    modport server (input  DDRARB, DMA0ACLK, DMA0DAREADY, DMA0DRLAST, DMA0DRTYPE, DMA0DRVALID, DMA1ACLK, DMA1DAREADY, DMA1DRLAST, DMA1DRTYPE, DMA1DRVALID, DMA2ACLK, DMA2DAREADY, DMA2DRLAST, DMA2DRTYPE, DMA2DRVALID, DMA3ACLK, DMA3DAREADY, DMA3DRLAST, DMA3DRTYPE, DMA3DRVALID, EMIOCAN0PHYRX, EMIOCAN1PHYRX, EMIOENET0EXTINTIN, EMIOENET0GMIICOL, EMIOENET0GMIICRS, EMIOENET0GMIIRXCLK, EMIOENET0GMIIRXD, EMIOENET0GMIIRXDV, EMIOENET0GMIIRXER, EMIOENET0GMIITXCLK, EMIOENET0MDIOI, EMIOENET1EXTINTIN, EMIOENET1GMIICOL, EMIOENET1GMIICRS, EMIOENET1GMIIRXCLK, EMIOENET1GMIIRXD, EMIOENET1GMIIRXDV, EMIOENET1GMIIRXER, EMIOENET1GMIITXCLK, EMIOENET1MDIOI, EMIOGPIOI, EMIOI2C0SCLI, EMIOI2C0SDAI, EMIOI2C1SCLI, EMIOI2C1SDAI, EMIOPJTAGTCK, EMIOPJTAGTDI, EMIOPJTAGTMS, EMIOSDIO0CDN, EMIOSDIO0CLKFB, EMIOSDIO0CMDI, EMIOSDIO0DATAI, EMIOSDIO0WP, EMIOSDIO1CDN, EMIOSDIO1CLKFB, EMIOSDIO1CMDI, EMIOSDIO1DATAI, EMIOSDIO1WP, EMIOSPI0MI, EMIOSPI0SCLKI, EMIOSPI0SI, EMIOSPI0SSIN, EMIOSPI1MI, EMIOSPI1SCLKI, EMIOSPI1SI, EMIOSPI1SSIN, EMIOSRAMINTIN, EMIOTRACECLK, EMIOTTC0CLKI, EMIOTTC1CLKI, EMIOUART0CTSN, EMIOUART0DCDN, EMIOUART0DSRN, EMIOUART0RIN, EMIOUART0RX, EMIOUART1CTSN, EMIOUART1DCDN, EMIOUART1DSRN, EMIOUART1RIN, EMIOUART1RX, EMIOUSB0VBUSPWRFAULT, EMIOUSB1VBUSPWRFAULT, EMIOWDTCLKI, EVENTEVENTI, FCLKCLKTRIGN, FPGAIDLEN, FTMDTRACEINATID, FTMDTRACEINCLOCK, FTMDTRACEINDATA, FTMDTRACEINVALID, FTMTF2PDEBUG, FTMTF2PTRIG, FTMTP2FTRIGACK, IRQF2P, MAXIGP0ACLK, MAXIGP0ARREADY, MAXIGP0AWREADY, MAXIGP0BID, MAXIGP0BRESP, MAXIGP0BVALID, MAXIGP0RDATA, MAXIGP0RID, MAXIGP0RLAST, MAXIGP0RRESP, MAXIGP0RVALID, MAXIGP0WREADY, MAXIGP1ACLK, MAXIGP1ARREADY, MAXIGP1AWREADY, MAXIGP1BID, MAXIGP1BRESP, MAXIGP1BVALID, MAXIGP1RDATA, MAXIGP1RID, MAXIGP1RLAST, MAXIGP1RRESP, MAXIGP1RVALID, MAXIGP1WREADY, SAXIACPACLK, SAXIACPARADDR, SAXIACPARBURST, SAXIACPARCACHE, SAXIACPARID, SAXIACPARLEN, SAXIACPARLOCK, SAXIACPARPROT, SAXIACPARQOS, SAXIACPARSIZE, SAXIACPARUSER, SAXIACPARVALID, SAXIACPAWADDR, SAXIACPAWBURST, SAXIACPAWCACHE, SAXIACPAWID, SAXIACPAWLEN, SAXIACPAWLOCK, SAXIACPAWPROT, SAXIACPAWQOS, SAXIACPAWSIZE, SAXIACPAWUSER, SAXIACPAWVALID, SAXIACPBREADY, SAXIACPRREADY, SAXIACPWDATA, SAXIACPWID, SAXIACPWLAST, SAXIACPWSTRB, SAXIACPWVALID, SAXIGP0ACLK, SAXIGP0ARADDR, SAXIGP0ARBURST, SAXIGP0ARCACHE, SAXIGP0ARID, SAXIGP0ARLEN, SAXIGP0ARLOCK, SAXIGP0ARPROT, SAXIGP0ARQOS, SAXIGP0ARSIZE, SAXIGP0ARVALID, SAXIGP0AWADDR, SAXIGP0AWBURST, SAXIGP0AWCACHE, SAXIGP0AWID, SAXIGP0AWLEN, SAXIGP0AWLOCK, SAXIGP0AWPROT, SAXIGP0AWQOS, SAXIGP0AWSIZE, SAXIGP0AWVALID, SAXIGP0BREADY, SAXIGP0RREADY, SAXIGP0WDATA, SAXIGP0WID, SAXIGP0WLAST, SAXIGP0WSTRB, SAXIGP0WVALID, SAXIGP1ACLK, SAXIGP1ARADDR, SAXIGP1ARBURST, SAXIGP1ARCACHE, SAXIGP1ARID, SAXIGP1ARLEN, SAXIGP1ARLOCK, SAXIGP1ARPROT, SAXIGP1ARQOS, SAXIGP1ARSIZE, SAXIGP1ARVALID, SAXIGP1AWADDR, SAXIGP1AWBURST, SAXIGP1AWCACHE, SAXIGP1AWID, SAXIGP1AWLEN, SAXIGP1AWLOCK, SAXIGP1AWPROT, SAXIGP1AWQOS, SAXIGP1AWSIZE, SAXIGP1AWVALID, SAXIGP1BREADY, SAXIGP1RREADY, SAXIGP1WDATA, SAXIGP1WID, SAXIGP1WLAST, SAXIGP1WSTRB, SAXIGP1WVALID, SAXIHP0ACLK, SAXIHP0ARADDR, SAXIHP0ARBURST, SAXIHP0ARCACHE, SAXIHP0ARID, SAXIHP0ARLEN, SAXIHP0ARLOCK, SAXIHP0ARPROT, SAXIHP0ARQOS, SAXIHP0ARSIZE, SAXIHP0ARVALID, SAXIHP0AWADDR, SAXIHP0AWBURST, SAXIHP0AWCACHE, SAXIHP0AWID, SAXIHP0AWLEN, SAXIHP0AWLOCK, SAXIHP0AWPROT, SAXIHP0AWQOS, SAXIHP0AWSIZE, SAXIHP0AWVALID, SAXIHP0BREADY, SAXIHP0RDISSUECAP1EN, SAXIHP0RREADY, SAXIHP0WDATA, SAXIHP0WID, SAXIHP0WLAST, SAXIHP0WRISSUECAP1EN, SAXIHP0WSTRB, SAXIHP0WVALID, SAXIHP1ACLK, SAXIHP1ARADDR, SAXIHP1ARBURST, SAXIHP1ARCACHE, SAXIHP1ARID, SAXIHP1ARLEN, SAXIHP1ARLOCK, SAXIHP1ARPROT, SAXIHP1ARQOS, SAXIHP1ARSIZE, SAXIHP1ARVALID, SAXIHP1AWADDR, SAXIHP1AWBURST, SAXIHP1AWCACHE, SAXIHP1AWID, SAXIHP1AWLEN, SAXIHP1AWLOCK, SAXIHP1AWPROT, SAXIHP1AWQOS, SAXIHP1AWSIZE, SAXIHP1AWVALID, SAXIHP1BREADY, SAXIHP1RDISSUECAP1EN, SAXIHP1RREADY, SAXIHP1WDATA, SAXIHP1WID, SAXIHP1WLAST, SAXIHP1WRISSUECAP1EN, SAXIHP1WSTRB, SAXIHP1WVALID, SAXIHP2ACLK, SAXIHP2ARADDR, SAXIHP2ARBURST, SAXIHP2ARCACHE, SAXIHP2ARID, SAXIHP2ARLEN, SAXIHP2ARLOCK, SAXIHP2ARPROT, SAXIHP2ARQOS, SAXIHP2ARSIZE, SAXIHP2ARVALID, SAXIHP2AWADDR, SAXIHP2AWBURST, SAXIHP2AWCACHE, SAXIHP2AWID, SAXIHP2AWLEN, SAXIHP2AWLOCK, SAXIHP2AWPROT, SAXIHP2AWQOS, SAXIHP2AWSIZE, SAXIHP2AWVALID, SAXIHP2BREADY, SAXIHP2RDISSUECAP1EN, SAXIHP2RREADY, SAXIHP2WDATA, SAXIHP2WID, SAXIHP2WLAST, SAXIHP2WRISSUECAP1EN, SAXIHP2WSTRB, SAXIHP2WVALID, SAXIHP3ACLK, SAXIHP3ARADDR, SAXIHP3ARBURST, SAXIHP3ARCACHE, SAXIHP3ARID, SAXIHP3ARLEN, SAXIHP3ARLOCK, SAXIHP3ARPROT, SAXIHP3ARQOS, SAXIHP3ARSIZE, SAXIHP3ARVALID, SAXIHP3AWADDR, SAXIHP3AWBURST, SAXIHP3AWCACHE, SAXIHP3AWID, SAXIHP3AWLEN, SAXIHP3AWLOCK, SAXIHP3AWPROT, SAXIHP3AWQOS, SAXIHP3AWSIZE, SAXIHP3AWVALID, SAXIHP3BREADY, SAXIHP3RDISSUECAP1EN, SAXIHP3RREADY, SAXIHP3WDATA, SAXIHP3WID, SAXIHP3WLAST, SAXIHP3WRISSUECAP1EN, SAXIHP3WSTRB, SAXIHP3WVALID,
                    output DMA0DATYPE, DMA0DAVALID, DMA0DRREADY, DMA0RSTN, DMA1DATYPE, DMA1DAVALID, DMA1DRREADY, DMA1RSTN, DMA2DATYPE, DMA2DAVALID, DMA2DRREADY, DMA2RSTN, DMA3DATYPE, DMA3DAVALID, DMA3DRREADY, DMA3RSTN, EMIOCAN0PHYTX, EMIOCAN1PHYTX, EMIOENET0GMIITXD, EMIOENET0GMIITXEN, EMIOENET0GMIITXER, EMIOENET0MDIOMDC, EMIOENET0MDIOO, EMIOENET0MDIOTN, EMIOENET0PTPDELAYREQRX, EMIOENET0PTPDELAYREQTX, EMIOENET0PTPPDELAYREQRX, EMIOENET0PTPPDELAYREQTX, EMIOENET0PTPPDELAYRESPRX, EMIOENET0PTPPDELAYRESPTX, EMIOENET0PTPSYNCFRAMERX, EMIOENET0PTPSYNCFRAMETX, EMIOENET0SOFRX, EMIOENET0SOFTX, EMIOENET1GMIITXD, EMIOENET1GMIITXEN, EMIOENET1GMIITXER, EMIOENET1MDIOMDC, EMIOENET1MDIOO, EMIOENET1MDIOTN, EMIOENET1PTPDELAYREQRX, EMIOENET1PTPDELAYREQTX, EMIOENET1PTPPDELAYREQRX, EMIOENET1PTPPDELAYREQTX, EMIOENET1PTPPDELAYRESPRX, EMIOENET1PTPPDELAYRESPTX, EMIOENET1PTPSYNCFRAMERX, EMIOENET1PTPSYNCFRAMETX, EMIOENET1SOFRX, EMIOENET1SOFTX, EMIOGPIOO, EMIOGPIOTN, EMIOI2C0SCLO, EMIOI2C0SCLTN, EMIOI2C0SDAO, EMIOI2C0SDATN, EMIOI2C1SCLO, EMIOI2C1SCLTN, EMIOI2C1SDAO, EMIOI2C1SDATN, EMIOPJTAGTDO, EMIOPJTAGTDTN, EMIOSDIO0BUSPOW, EMIOSDIO0BUSVOLT, EMIOSDIO0CLK, EMIOSDIO0CMDO, EMIOSDIO0CMDTN, EMIOSDIO0DATAO, EMIOSDIO0DATATN, EMIOSDIO0LED, EMIOSDIO1BUSPOW, EMIOSDIO1BUSVOLT, EMIOSDIO1CLK, EMIOSDIO1CMDO, EMIOSDIO1CMDTN, EMIOSDIO1DATAO, EMIOSDIO1DATATN, EMIOSDIO1LED, EMIOSPI0MO, EMIOSPI0MOTN, EMIOSPI0SCLKO, EMIOSPI0SCLKTN, EMIOSPI0SO, EMIOSPI0SSNTN, EMIOSPI0SSON, EMIOSPI0STN, EMIOSPI1MO, EMIOSPI1MOTN, EMIOSPI1SCLKO, EMIOSPI1SCLKTN, EMIOSPI1SO, EMIOSPI1SSNTN, EMIOSPI1SSON, EMIOSPI1STN, EMIOTRACECTL, EMIOTRACEDATA, EMIOTTC0WAVEO, EMIOTTC1WAVEO, EMIOUART0DTRN, EMIOUART0RTSN, EMIOUART0TX, EMIOUART1DTRN, EMIOUART1RTSN, EMIOUART1TX, EMIOUSB0PORTINDCTL, EMIOUSB0VBUSPWRSELECT, EMIOUSB1PORTINDCTL, EMIOUSB1VBUSPWRSELECT, EMIOWDTRSTO, EVENTEVENTO, EVENTSTANDBYWFE, EVENTSTANDBYWFI, FCLKCLK, FCLKRESETN, FTMTF2PTRIGACK, FTMTP2FDEBUG, FTMTP2FTRIG, IRQP2F, MAXIGP0ARADDR, MAXIGP0ARBURST, MAXIGP0ARCACHE, MAXIGP0ARESETN, MAXIGP0ARID, MAXIGP0ARLEN, MAXIGP0ARLOCK, MAXIGP0ARPROT, MAXIGP0ARQOS, MAXIGP0ARSIZE, MAXIGP0ARVALID, MAXIGP0AWADDR, MAXIGP0AWBURST, MAXIGP0AWCACHE, MAXIGP0AWID, MAXIGP0AWLEN, MAXIGP0AWLOCK, MAXIGP0AWPROT, MAXIGP0AWQOS, MAXIGP0AWSIZE, MAXIGP0AWVALID, MAXIGP0BREADY, MAXIGP0RREADY, MAXIGP0WDATA, MAXIGP0WID, MAXIGP0WLAST, MAXIGP0WSTRB, MAXIGP0WVALID, MAXIGP1ARADDR, MAXIGP1ARBURST, MAXIGP1ARCACHE, MAXIGP1ARESETN, MAXIGP1ARID, MAXIGP1ARLEN, MAXIGP1ARLOCK, MAXIGP1ARPROT, MAXIGP1ARQOS, MAXIGP1ARSIZE, MAXIGP1ARVALID, MAXIGP1AWADDR, MAXIGP1AWBURST, MAXIGP1AWCACHE, MAXIGP1AWID, MAXIGP1AWLEN, MAXIGP1AWLOCK, MAXIGP1AWPROT, MAXIGP1AWQOS, MAXIGP1AWSIZE, MAXIGP1AWVALID, MAXIGP1BREADY, MAXIGP1RREADY, MAXIGP1WDATA, MAXIGP1WID, MAXIGP1WLAST, MAXIGP1WSTRB, MAXIGP1WVALID, SAXIACPARESETN, SAXIACPARREADY, SAXIACPAWREADY, SAXIACPBID, SAXIACPBRESP, SAXIACPBVALID, SAXIACPRDATA, SAXIACPRID, SAXIACPRLAST, SAXIACPRRESP, SAXIACPRVALID, SAXIACPWREADY, SAXIGP0ARESETN, SAXIGP0ARREADY, SAXIGP0AWREADY, SAXIGP0BID, SAXIGP0BRESP, SAXIGP0BVALID, SAXIGP0RDATA, SAXIGP0RID, SAXIGP0RLAST, SAXIGP0RRESP, SAXIGP0RVALID, SAXIGP0WREADY, SAXIGP1ARESETN, SAXIGP1ARREADY, SAXIGP1AWREADY, SAXIGP1BID, SAXIGP1BRESP, SAXIGP1BVALID, SAXIGP1RDATA, SAXIGP1RID, SAXIGP1RLAST, SAXIGP1RRESP, SAXIGP1RVALID, SAXIGP1WREADY, SAXIHP0ARESETN, SAXIHP0ARREADY, SAXIHP0AWREADY, SAXIHP0BID, SAXIHP0BRESP, SAXIHP0BVALID, SAXIHP0RACOUNT, SAXIHP0RCOUNT, SAXIHP0RDATA, SAXIHP0RID, SAXIHP0RLAST, SAXIHP0RRESP, SAXIHP0RVALID, SAXIHP0WACOUNT, SAXIHP0WCOUNT, SAXIHP0WREADY, SAXIHP1ARESETN, SAXIHP1ARREADY, SAXIHP1AWREADY, SAXIHP1BID, SAXIHP1BRESP, SAXIHP1BVALID, SAXIHP1RACOUNT, SAXIHP1RCOUNT, SAXIHP1RDATA, SAXIHP1RID, SAXIHP1RLAST, SAXIHP1RRESP, SAXIHP1RVALID, SAXIHP1WACOUNT, SAXIHP1WCOUNT, SAXIHP1WREADY, SAXIHP2ARESETN, SAXIHP2ARREADY, SAXIHP2AWREADY, SAXIHP2BID, SAXIHP2BRESP, SAXIHP2BVALID, SAXIHP2RACOUNT, SAXIHP2RCOUNT, SAXIHP2RDATA, SAXIHP2RID, SAXIHP2RLAST, SAXIHP2RRESP, SAXIHP2RVALID, SAXIHP2WACOUNT, SAXIHP2WCOUNT, SAXIHP2WREADY, SAXIHP3ARESETN, SAXIHP3ARREADY, SAXIHP3AWREADY, SAXIHP3BID, SAXIHP3BRESP, SAXIHP3BVALID, SAXIHP3RACOUNT, SAXIHP3RCOUNT, SAXIHP3RDATA, SAXIHP3RID, SAXIHP3RLAST, SAXIHP3RRESP, SAXIHP3RVALID, SAXIHP3WACOUNT, SAXIHP3WCOUNT, SAXIHP3WREADY);
    modport client (output DDRARB, DMA0ACLK, DMA0DAREADY, DMA0DRLAST, DMA0DRTYPE, DMA0DRVALID, DMA1ACLK, DMA1DAREADY, DMA1DRLAST, DMA1DRTYPE, DMA1DRVALID, DMA2ACLK, DMA2DAREADY, DMA2DRLAST, DMA2DRTYPE, DMA2DRVALID, DMA3ACLK, DMA3DAREADY, DMA3DRLAST, DMA3DRTYPE, DMA3DRVALID, EMIOCAN0PHYRX, EMIOCAN1PHYRX, EMIOENET0EXTINTIN, EMIOENET0GMIICOL, EMIOENET0GMIICRS, EMIOENET0GMIIRXCLK, EMIOENET0GMIIRXD, EMIOENET0GMIIRXDV, EMIOENET0GMIIRXER, EMIOENET0GMIITXCLK, EMIOENET0MDIOI, EMIOENET1EXTINTIN, EMIOENET1GMIICOL, EMIOENET1GMIICRS, EMIOENET1GMIIRXCLK, EMIOENET1GMIIRXD, EMIOENET1GMIIRXDV, EMIOENET1GMIIRXER, EMIOENET1GMIITXCLK, EMIOENET1MDIOI, EMIOGPIOI, EMIOI2C0SCLI, EMIOI2C0SDAI, EMIOI2C1SCLI, EMIOI2C1SDAI, EMIOPJTAGTCK, EMIOPJTAGTDI, EMIOPJTAGTMS, EMIOSDIO0CDN, EMIOSDIO0CLKFB, EMIOSDIO0CMDI, EMIOSDIO0DATAI, EMIOSDIO0WP, EMIOSDIO1CDN, EMIOSDIO1CLKFB, EMIOSDIO1CMDI, EMIOSDIO1DATAI, EMIOSDIO1WP, EMIOSPI0MI, EMIOSPI0SCLKI, EMIOSPI0SI, EMIOSPI0SSIN, EMIOSPI1MI, EMIOSPI1SCLKI, EMIOSPI1SI, EMIOSPI1SSIN, EMIOSRAMINTIN, EMIOTRACECLK, EMIOTTC0CLKI, EMIOTTC1CLKI, EMIOUART0CTSN, EMIOUART0DCDN, EMIOUART0DSRN, EMIOUART0RIN, EMIOUART0RX, EMIOUART1CTSN, EMIOUART1DCDN, EMIOUART1DSRN, EMIOUART1RIN, EMIOUART1RX, EMIOUSB0VBUSPWRFAULT, EMIOUSB1VBUSPWRFAULT, EMIOWDTCLKI, EVENTEVENTI, FCLKCLKTRIGN, FPGAIDLEN, FTMDTRACEINATID, FTMDTRACEINCLOCK, FTMDTRACEINDATA, FTMDTRACEINVALID, FTMTF2PDEBUG, FTMTF2PTRIG, FTMTP2FTRIGACK, IRQF2P, MAXIGP0ACLK, MAXIGP0ARREADY, MAXIGP0AWREADY, MAXIGP0BID, MAXIGP0BRESP, MAXIGP0BVALID, MAXIGP0RDATA, MAXIGP0RID, MAXIGP0RLAST, MAXIGP0RRESP, MAXIGP0RVALID, MAXIGP0WREADY, MAXIGP1ACLK, MAXIGP1ARREADY, MAXIGP1AWREADY, MAXIGP1BID, MAXIGP1BRESP, MAXIGP1BVALID, MAXIGP1RDATA, MAXIGP1RID, MAXIGP1RLAST, MAXIGP1RRESP, MAXIGP1RVALID, MAXIGP1WREADY, SAXIACPACLK, SAXIACPARADDR, SAXIACPARBURST, SAXIACPARCACHE, SAXIACPARID, SAXIACPARLEN, SAXIACPARLOCK, SAXIACPARPROT, SAXIACPARQOS, SAXIACPARSIZE, SAXIACPARUSER, SAXIACPARVALID, SAXIACPAWADDR, SAXIACPAWBURST, SAXIACPAWCACHE, SAXIACPAWID, SAXIACPAWLEN, SAXIACPAWLOCK, SAXIACPAWPROT, SAXIACPAWQOS, SAXIACPAWSIZE, SAXIACPAWUSER, SAXIACPAWVALID, SAXIACPBREADY, SAXIACPRREADY, SAXIACPWDATA, SAXIACPWID, SAXIACPWLAST, SAXIACPWSTRB, SAXIACPWVALID, SAXIGP0ACLK, SAXIGP0ARADDR, SAXIGP0ARBURST, SAXIGP0ARCACHE, SAXIGP0ARID, SAXIGP0ARLEN, SAXIGP0ARLOCK, SAXIGP0ARPROT, SAXIGP0ARQOS, SAXIGP0ARSIZE, SAXIGP0ARVALID, SAXIGP0AWADDR, SAXIGP0AWBURST, SAXIGP0AWCACHE, SAXIGP0AWID, SAXIGP0AWLEN, SAXIGP0AWLOCK, SAXIGP0AWPROT, SAXIGP0AWQOS, SAXIGP0AWSIZE, SAXIGP0AWVALID, SAXIGP0BREADY, SAXIGP0RREADY, SAXIGP0WDATA, SAXIGP0WID, SAXIGP0WLAST, SAXIGP0WSTRB, SAXIGP0WVALID, SAXIGP1ACLK, SAXIGP1ARADDR, SAXIGP1ARBURST, SAXIGP1ARCACHE, SAXIGP1ARID, SAXIGP1ARLEN, SAXIGP1ARLOCK, SAXIGP1ARPROT, SAXIGP1ARQOS, SAXIGP1ARSIZE, SAXIGP1ARVALID, SAXIGP1AWADDR, SAXIGP1AWBURST, SAXIGP1AWCACHE, SAXIGP1AWID, SAXIGP1AWLEN, SAXIGP1AWLOCK, SAXIGP1AWPROT, SAXIGP1AWQOS, SAXIGP1AWSIZE, SAXIGP1AWVALID, SAXIGP1BREADY, SAXIGP1RREADY, SAXIGP1WDATA, SAXIGP1WID, SAXIGP1WLAST, SAXIGP1WSTRB, SAXIGP1WVALID, SAXIHP0ACLK, SAXIHP0ARADDR, SAXIHP0ARBURST, SAXIHP0ARCACHE, SAXIHP0ARID, SAXIHP0ARLEN, SAXIHP0ARLOCK, SAXIHP0ARPROT, SAXIHP0ARQOS, SAXIHP0ARSIZE, SAXIHP0ARVALID, SAXIHP0AWADDR, SAXIHP0AWBURST, SAXIHP0AWCACHE, SAXIHP0AWID, SAXIHP0AWLEN, SAXIHP0AWLOCK, SAXIHP0AWPROT, SAXIHP0AWQOS, SAXIHP0AWSIZE, SAXIHP0AWVALID, SAXIHP0BREADY, SAXIHP0RDISSUECAP1EN, SAXIHP0RREADY, SAXIHP0WDATA, SAXIHP0WID, SAXIHP0WLAST, SAXIHP0WRISSUECAP1EN, SAXIHP0WSTRB, SAXIHP0WVALID, SAXIHP1ACLK, SAXIHP1ARADDR, SAXIHP1ARBURST, SAXIHP1ARCACHE, SAXIHP1ARID, SAXIHP1ARLEN, SAXIHP1ARLOCK, SAXIHP1ARPROT, SAXIHP1ARQOS, SAXIHP1ARSIZE, SAXIHP1ARVALID, SAXIHP1AWADDR, SAXIHP1AWBURST, SAXIHP1AWCACHE, SAXIHP1AWID, SAXIHP1AWLEN, SAXIHP1AWLOCK, SAXIHP1AWPROT, SAXIHP1AWQOS, SAXIHP1AWSIZE, SAXIHP1AWVALID, SAXIHP1BREADY, SAXIHP1RDISSUECAP1EN, SAXIHP1RREADY, SAXIHP1WDATA, SAXIHP1WID, SAXIHP1WLAST, SAXIHP1WRISSUECAP1EN, SAXIHP1WSTRB, SAXIHP1WVALID, SAXIHP2ACLK, SAXIHP2ARADDR, SAXIHP2ARBURST, SAXIHP2ARCACHE, SAXIHP2ARID, SAXIHP2ARLEN, SAXIHP2ARLOCK, SAXIHP2ARPROT, SAXIHP2ARQOS, SAXIHP2ARSIZE, SAXIHP2ARVALID, SAXIHP2AWADDR, SAXIHP2AWBURST, SAXIHP2AWCACHE, SAXIHP2AWID, SAXIHP2AWLEN, SAXIHP2AWLOCK, SAXIHP2AWPROT, SAXIHP2AWQOS, SAXIHP2AWSIZE, SAXIHP2AWVALID, SAXIHP2BREADY, SAXIHP2RDISSUECAP1EN, SAXIHP2RREADY, SAXIHP2WDATA, SAXIHP2WID, SAXIHP2WLAST, SAXIHP2WRISSUECAP1EN, SAXIHP2WSTRB, SAXIHP2WVALID, SAXIHP3ACLK, SAXIHP3ARADDR, SAXIHP3ARBURST, SAXIHP3ARCACHE, SAXIHP3ARID, SAXIHP3ARLEN, SAXIHP3ARLOCK, SAXIHP3ARPROT, SAXIHP3ARQOS, SAXIHP3ARSIZE, SAXIHP3ARVALID, SAXIHP3AWADDR, SAXIHP3AWBURST, SAXIHP3AWCACHE, SAXIHP3AWID, SAXIHP3AWLEN, SAXIHP3AWLOCK, SAXIHP3AWPROT, SAXIHP3AWQOS, SAXIHP3AWSIZE, SAXIHP3AWVALID, SAXIHP3BREADY, SAXIHP3RDISSUECAP1EN, SAXIHP3RREADY, SAXIHP3WDATA, SAXIHP3WID, SAXIHP3WLAST, SAXIHP3WRISSUECAP1EN, SAXIHP3WSTRB, SAXIHP3WVALID,
                    input  DMA0DATYPE, DMA0DAVALID, DMA0DRREADY, DMA0RSTN, DMA1DATYPE, DMA1DAVALID, DMA1DRREADY, DMA1RSTN, DMA2DATYPE, DMA2DAVALID, DMA2DRREADY, DMA2RSTN, DMA3DATYPE, DMA3DAVALID, DMA3DRREADY, DMA3RSTN, EMIOCAN0PHYTX, EMIOCAN1PHYTX, EMIOENET0GMIITXD, EMIOENET0GMIITXEN, EMIOENET0GMIITXER, EMIOENET0MDIOMDC, EMIOENET0MDIOO, EMIOENET0MDIOTN, EMIOENET0PTPDELAYREQRX, EMIOENET0PTPDELAYREQTX, EMIOENET0PTPPDELAYREQRX, EMIOENET0PTPPDELAYREQTX, EMIOENET0PTPPDELAYRESPRX, EMIOENET0PTPPDELAYRESPTX, EMIOENET0PTPSYNCFRAMERX, EMIOENET0PTPSYNCFRAMETX, EMIOENET0SOFRX, EMIOENET0SOFTX, EMIOENET1GMIITXD, EMIOENET1GMIITXEN, EMIOENET1GMIITXER, EMIOENET1MDIOMDC, EMIOENET1MDIOO, EMIOENET1MDIOTN, EMIOENET1PTPDELAYREQRX, EMIOENET1PTPDELAYREQTX, EMIOENET1PTPPDELAYREQRX, EMIOENET1PTPPDELAYREQTX, EMIOENET1PTPPDELAYRESPRX, EMIOENET1PTPPDELAYRESPTX, EMIOENET1PTPSYNCFRAMERX, EMIOENET1PTPSYNCFRAMETX, EMIOENET1SOFRX, EMIOENET1SOFTX, EMIOGPIOO, EMIOGPIOTN, EMIOI2C0SCLO, EMIOI2C0SCLTN, EMIOI2C0SDAO, EMIOI2C0SDATN, EMIOI2C1SCLO, EMIOI2C1SCLTN, EMIOI2C1SDAO, EMIOI2C1SDATN, EMIOPJTAGTDO, EMIOPJTAGTDTN, EMIOSDIO0BUSPOW, EMIOSDIO0BUSVOLT, EMIOSDIO0CLK, EMIOSDIO0CMDO, EMIOSDIO0CMDTN, EMIOSDIO0DATAO, EMIOSDIO0DATATN, EMIOSDIO0LED, EMIOSDIO1BUSPOW, EMIOSDIO1BUSVOLT, EMIOSDIO1CLK, EMIOSDIO1CMDO, EMIOSDIO1CMDTN, EMIOSDIO1DATAO, EMIOSDIO1DATATN, EMIOSDIO1LED, EMIOSPI0MO, EMIOSPI0MOTN, EMIOSPI0SCLKO, EMIOSPI0SCLKTN, EMIOSPI0SO, EMIOSPI0SSNTN, EMIOSPI0SSON, EMIOSPI0STN, EMIOSPI1MO, EMIOSPI1MOTN, EMIOSPI1SCLKO, EMIOSPI1SCLKTN, EMIOSPI1SO, EMIOSPI1SSNTN, EMIOSPI1SSON, EMIOSPI1STN, EMIOTRACECTL, EMIOTRACEDATA, EMIOTTC0WAVEO, EMIOTTC1WAVEO, EMIOUART0DTRN, EMIOUART0RTSN, EMIOUART0TX, EMIOUART1DTRN, EMIOUART1RTSN, EMIOUART1TX, EMIOUSB0PORTINDCTL, EMIOUSB0VBUSPWRSELECT, EMIOUSB1PORTINDCTL, EMIOUSB1VBUSPWRSELECT, EMIOWDTRSTO, EVENTEVENTO, EVENTSTANDBYWFE, EVENTSTANDBYWFI, FCLKCLK, FCLKRESETN, FTMTF2PTRIGACK, FTMTP2FDEBUG, FTMTP2FTRIG, IRQP2F, MAXIGP0ARADDR, MAXIGP0ARBURST, MAXIGP0ARCACHE, MAXIGP0ARESETN, MAXIGP0ARID, MAXIGP0ARLEN, MAXIGP0ARLOCK, MAXIGP0ARPROT, MAXIGP0ARQOS, MAXIGP0ARSIZE, MAXIGP0ARVALID, MAXIGP0AWADDR, MAXIGP0AWBURST, MAXIGP0AWCACHE, MAXIGP0AWID, MAXIGP0AWLEN, MAXIGP0AWLOCK, MAXIGP0AWPROT, MAXIGP0AWQOS, MAXIGP0AWSIZE, MAXIGP0AWVALID, MAXIGP0BREADY, MAXIGP0RREADY, MAXIGP0WDATA, MAXIGP0WID, MAXIGP0WLAST, MAXIGP0WSTRB, MAXIGP0WVALID, MAXIGP1ARADDR, MAXIGP1ARBURST, MAXIGP1ARCACHE, MAXIGP1ARESETN, MAXIGP1ARID, MAXIGP1ARLEN, MAXIGP1ARLOCK, MAXIGP1ARPROT, MAXIGP1ARQOS, MAXIGP1ARSIZE, MAXIGP1ARVALID, MAXIGP1AWADDR, MAXIGP1AWBURST, MAXIGP1AWCACHE, MAXIGP1AWID, MAXIGP1AWLEN, MAXIGP1AWLOCK, MAXIGP1AWPROT, MAXIGP1AWQOS, MAXIGP1AWSIZE, MAXIGP1AWVALID, MAXIGP1BREADY, MAXIGP1RREADY, MAXIGP1WDATA, MAXIGP1WID, MAXIGP1WLAST, MAXIGP1WSTRB, MAXIGP1WVALID, SAXIACPARESETN, SAXIACPARREADY, SAXIACPAWREADY, SAXIACPBID, SAXIACPBRESP, SAXIACPBVALID, SAXIACPRDATA, SAXIACPRID, SAXIACPRLAST, SAXIACPRRESP, SAXIACPRVALID, SAXIACPWREADY, SAXIGP0ARESETN, SAXIGP0ARREADY, SAXIGP0AWREADY, SAXIGP0BID, SAXIGP0BRESP, SAXIGP0BVALID, SAXIGP0RDATA, SAXIGP0RID, SAXIGP0RLAST, SAXIGP0RRESP, SAXIGP0RVALID, SAXIGP0WREADY, SAXIGP1ARESETN, SAXIGP1ARREADY, SAXIGP1AWREADY, SAXIGP1BID, SAXIGP1BRESP, SAXIGP1BVALID, SAXIGP1RDATA, SAXIGP1RID, SAXIGP1RLAST, SAXIGP1RRESP, SAXIGP1RVALID, SAXIGP1WREADY, SAXIHP0ARESETN, SAXIHP0ARREADY, SAXIHP0AWREADY, SAXIHP0BID, SAXIHP0BRESP, SAXIHP0BVALID, SAXIHP0RACOUNT, SAXIHP0RCOUNT, SAXIHP0RDATA, SAXIHP0RID, SAXIHP0RLAST, SAXIHP0RRESP, SAXIHP0RVALID, SAXIHP0WACOUNT, SAXIHP0WCOUNT, SAXIHP0WREADY, SAXIHP1ARESETN, SAXIHP1ARREADY, SAXIHP1AWREADY, SAXIHP1BID, SAXIHP1BRESP, SAXIHP1BVALID, SAXIHP1RACOUNT, SAXIHP1RCOUNT, SAXIHP1RDATA, SAXIHP1RID, SAXIHP1RLAST, SAXIHP1RRESP, SAXIHP1RVALID, SAXIHP1WACOUNT, SAXIHP1WCOUNT, SAXIHP1WREADY, SAXIHP2ARESETN, SAXIHP2ARREADY, SAXIHP2AWREADY, SAXIHP2BID, SAXIHP2BRESP, SAXIHP2BVALID, SAXIHP2RACOUNT, SAXIHP2RCOUNT, SAXIHP2RDATA, SAXIHP2RID, SAXIHP2RLAST, SAXIHP2RRESP, SAXIHP2RVALID, SAXIHP2WACOUNT, SAXIHP2WCOUNT, SAXIHP2WREADY, SAXIHP3ARESETN, SAXIHP3ARREADY, SAXIHP3AWREADY, SAXIHP3BID, SAXIHP3BRESP, SAXIHP3BVALID, SAXIHP3RACOUNT, SAXIHP3RCOUNT, SAXIHP3RDATA, SAXIHP3RID, SAXIHP3RLAST, SAXIHP3RRESP, SAXIHP3RVALID, SAXIHP3WACOUNT, SAXIHP3WCOUNT, SAXIHP3WREADY);
endinterface
`endif
`ifndef __ZynqTopIFC_DEF__
`define __ZynqTopIFC_DEF__
interface ZynqTopIFC;
    logic [54 - 1:0] MIO;
endinterface
`endif
//METASTART; P7Wrap
//METAINTERNAL; pps; PS7;
//METAINTERNAL; pclockTop; ClockTop;
//METAGUARD; MAXIGP0_I.R; 0 != pps$MAXIGP0RREADY;
//METAGUARD; MAXIGP0_I.B; 0 != pps$MAXIGP0BREADY;
//METAGUARD; RULE$init; 1;
//METAINVOKE; RULE$gp0ar__ENA; :MAXIGP0_O.AR__ENA;
//METAGUARD; RULE$gp0ar; !( ( 0 == pps$MAXIGP0ARVALID ) || ( !MAXIGP0_O.AR__RDY ) );
//METAINVOKE; RULE$gp0aw__ENA; :MAXIGP0_O.AW__ENA;
//METAGUARD; RULE$gp0aw; !( ( 0 == pps$MAXIGP0AWVALID ) || ( !MAXIGP0_O.AW__RDY ) );
//METAINVOKE; RULE$gp0w__ENA; :MAXIGP0_O.W__ENA;
//METAGUARD; RULE$gp0w; !( ( 0 == pps$MAXIGP0WVALID ) || ( !MAXIGP0_O.W__RDY ) );
//METARULES; RULE$init; RULE$gp0ar; RULE$gp0aw; RULE$gp0w
//METASTART; ZynqTop
//METAINTERNAL; ps7_ps7_foo; P7Wrap;
//METAINTERNAL; test; AxiTop;
//METAINTERNAL; ps7_fclk_0_c; BUFG;
//METAINTERNAL; ps7_freset_0_r; BUFG;
//METAGUARD; RULE$init; 1;
//METARULES; RULE$init
//METACONNECT; test$MAXIGP0_O.AR__ENA; ps7_ps7_foo$MAXIGP0_O.AR__ENA
//METACONNECT; test$MAXIGP0_O.AR__RDY; ps7_ps7_foo$MAXIGP0_O.AR__RDY
//METACONNECT; test$MAXIGP0_O.AW__ENA; ps7_ps7_foo$MAXIGP0_O.AW__ENA
//METACONNECT; test$MAXIGP0_O.AW__RDY; ps7_ps7_foo$MAXIGP0_O.AW__RDY
//METACONNECT; test$MAXIGP0_O.W__ENA; ps7_ps7_foo$MAXIGP0_O.W__ENA
//METACONNECT; test$MAXIGP0_O.W__RDY; ps7_ps7_foo$MAXIGP0_O.W__RDY
//METACONNECT; test$MAXIGP0_I.R__ENA; ps7_ps7_foo$MAXIGP0_I.R__ENA
//METACONNECT; test$MAXIGP0_I.R__RDY; ps7_ps7_foo$MAXIGP0_I.R__RDY
//METACONNECT; test$MAXIGP0_I.B__ENA; ps7_ps7_foo$MAXIGP0_I.B__ENA
//METACONNECT; test$MAXIGP0_I.B__RDY; ps7_ps7_foo$MAXIGP0_I.B__RDY
`endif
