`ifndef __fifo_GENERATED__VH__
`define __fifo_GENERATED__VH__

`endif
